module argTable(input clk, input [9:0] addr, output reg [15:0] data);
reg [15:0] mem [0:1023];
initial mem[0] = 16'h0;
initial mem[1] = 16'h3fff;
initial mem[2] = 16'h3fff;
initial mem[3] = 16'h3fff;
initial mem[4] = 16'h3fff;
initial mem[5] = 16'h3fff;
initial mem[6] = 16'h3fff;
initial mem[7] = 16'h3fff;
initial mem[8] = 16'h3fff;
initial mem[9] = 16'h3fff;
initial mem[10] = 16'h3fff;
initial mem[11] = 16'h3fff;
initial mem[12] = 16'h3fff;
initial mem[13] = 16'h3fff;
initial mem[14] = 16'h3fff;
initial mem[15] = 16'h3fff;
initial mem[16] = 16'hc001;
initial mem[17] = 16'hc001;
initial mem[18] = 16'hc001;
initial mem[19] = 16'hc001;
initial mem[20] = 16'hc001;
initial mem[21] = 16'hc001;
initial mem[22] = 16'hc001;
initial mem[23] = 16'hc001;
initial mem[24] = 16'hc001;
initial mem[25] = 16'hc001;
initial mem[26] = 16'hc001;
initial mem[27] = 16'hc001;
initial mem[28] = 16'hc001;
initial mem[29] = 16'hc001;
initial mem[30] = 16'hc001;
initial mem[31] = 16'hc001;
initial mem[32] = 16'h0;
initial mem[33] = 16'h1fff;
initial mem[34] = 16'h2d1b;
initial mem[35] = 16'h32e3;
initial mem[36] = 16'h3604;
initial mem[37] = 16'h37f4;
initial mem[38] = 16'h3944;
initial mem[39] = 16'h3a37;
initial mem[40] = 16'h3aee;
initial mem[41] = 16'h3b7d;
initial mem[42] = 16'h3bef;
initial mem[43] = 16'h3c4d;
initial mem[44] = 16'h3c9c;
initial mem[45] = 16'h3cde;
initial mem[46] = 16'h3d17;
initial mem[47] = 16'h3d49;
initial mem[48] = 16'hc28c;
initial mem[49] = 16'hc2b7;
initial mem[50] = 16'hc2e9;
initial mem[51] = 16'hc322;
initial mem[52] = 16'hc364;
initial mem[53] = 16'hc3b3;
initial mem[54] = 16'hc411;
initial mem[55] = 16'hc483;
initial mem[56] = 16'hc512;
initial mem[57] = 16'hc5c9;
initial mem[58] = 16'hc6bc;
initial mem[59] = 16'hc80c;
initial mem[60] = 16'hc9fc;
initial mem[61] = 16'hcd1d;
initial mem[62] = 16'hd2e5;
initial mem[63] = 16'he001;
initial mem[64] = 16'h0;
initial mem[65] = 16'h12e3;
initial mem[66] = 16'h1fff;
initial mem[67] = 16'h280a;
initial mem[68] = 16'h2d1b;
initial mem[69] = 16'h307e;
initial mem[70] = 16'h32e3;
initial mem[71] = 16'h34a8;
initial mem[72] = 16'h3604;
initial mem[73] = 16'h3716;
initial mem[74] = 16'h37f4;
initial mem[75] = 16'h38ab;
initial mem[76] = 16'h3944;
initial mem[77] = 16'h39c7;
initial mem[78] = 16'h3a37;
initial mem[79] = 16'h3a98;
initial mem[80] = 16'hc512;
initial mem[81] = 16'hc568;
initial mem[82] = 16'hc5c9;
initial mem[83] = 16'hc639;
initial mem[84] = 16'hc6bc;
initial mem[85] = 16'hc755;
initial mem[86] = 16'hc80c;
initial mem[87] = 16'hc8ea;
initial mem[88] = 16'hc9fc;
initial mem[89] = 16'hcb58;
initial mem[90] = 16'hcd1d;
initial mem[91] = 16'hcf82;
initial mem[92] = 16'hd2e5;
initial mem[93] = 16'hd7f6;
initial mem[94] = 16'he001;
initial mem[95] = 16'hed1d;
initial mem[96] = 16'h0;
initial mem[97] = 16'hd1b;
initial mem[98] = 16'h17f4;
initial mem[99] = 16'h1fff;
initial mem[100] = 16'h25c7;
initial mem[101] = 16'h29fa;
initial mem[102] = 16'h2d1b;
initial mem[103] = 16'h2f80;
initial mem[104] = 16'h3161;
initial mem[105] = 16'h32e3;
initial mem[106] = 16'h341f;
initial mem[107] = 16'h3526;
initial mem[108] = 16'h3604;
initial mem[109] = 16'h36c1;
initial mem[110] = 16'h3765;
initial mem[111] = 16'h37f4;
initial mem[112] = 16'hc78e;
initial mem[113] = 16'hc80c;
initial mem[114] = 16'hc89b;
initial mem[115] = 16'hc93f;
initial mem[116] = 16'hc9fc;
initial mem[117] = 16'hcada;
initial mem[118] = 16'hcbe1;
initial mem[119] = 16'hcd1d;
initial mem[120] = 16'hce9f;
initial mem[121] = 16'hd080;
initial mem[122] = 16'hd2e5;
initial mem[123] = 16'hd606;
initial mem[124] = 16'hda39;
initial mem[125] = 16'he001;
initial mem[126] = 16'he80c;
initial mem[127] = 16'hf2e5;
initial mem[128] = 16'h0;
initial mem[129] = 16'h9fb;
initial mem[130] = 16'h12e3;
initial mem[131] = 16'h1a37;
initial mem[132] = 16'h1fff;
initial mem[133] = 16'h2481;
initial mem[134] = 16'h280a;
initial mem[135] = 16'h2ad8;
initial mem[136] = 16'h2d1b;
initial mem[137] = 16'h2ef5;
initial mem[138] = 16'h307e;
initial mem[139] = 16'h31c9;
initial mem[140] = 16'h32e3;
initial mem[141] = 16'h33d6;
initial mem[142] = 16'h34a8;
initial mem[143] = 16'h3561;
initial mem[144] = 16'hc9fc;
initial mem[145] = 16'hca9f;
initial mem[146] = 16'hcb58;
initial mem[147] = 16'hcc2a;
initial mem[148] = 16'hcd1d;
initial mem[149] = 16'hce37;
initial mem[150] = 16'hcf82;
initial mem[151] = 16'hd10b;
initial mem[152] = 16'hd2e5;
initial mem[153] = 16'hd528;
initial mem[154] = 16'hd7f6;
initial mem[155] = 16'hdb7f;
initial mem[156] = 16'he001;
initial mem[157] = 16'he5c9;
initial mem[158] = 16'hed1d;
initial mem[159] = 16'hf605;
initial mem[160] = 16'h0;
initial mem[161] = 16'h80a;
initial mem[162] = 16'hf80;
initial mem[163] = 16'h1604;
initial mem[164] = 16'h1b7d;
initial mem[165] = 16'h1fff;
initial mem[166] = 16'h23b1;
initial mem[167] = 16'h26ba;
initial mem[168] = 16'h293d;
initial mem[169] = 16'h2b56;
initial mem[170] = 16'h2d1b;
initial mem[171] = 16'h2e9d;
initial mem[172] = 16'h2fe9;
initial mem[173] = 16'h3109;
initial mem[174] = 16'h3205;
initial mem[175] = 16'h32e3;
initial mem[176] = 16'hcc58;
initial mem[177] = 16'hcd1d;
initial mem[178] = 16'hcdfb;
initial mem[179] = 16'hcef7;
initial mem[180] = 16'hd017;
initial mem[181] = 16'hd163;
initial mem[182] = 16'hd2e5;
initial mem[183] = 16'hd4aa;
initial mem[184] = 16'hd6c3;
initial mem[185] = 16'hd946;
initial mem[186] = 16'hdc4f;
initial mem[187] = 16'he001;
initial mem[188] = 16'he483;
initial mem[189] = 16'he9fc;
initial mem[190] = 16'hf080;
initial mem[191] = 16'hf7f6;
initial mem[192] = 16'h0;
initial mem[193] = 16'h6ba;
initial mem[194] = 16'hd1b;
initial mem[195] = 16'h12e3;
initial mem[196] = 16'h17f4;
initial mem[197] = 16'h1c4e;
initial mem[198] = 16'h1fff;
initial mem[199] = 16'h2320;
initial mem[200] = 16'h25c7;
initial mem[201] = 16'h280a;
initial mem[202] = 16'h29fa;
initial mem[203] = 16'h2ba7;
initial mem[204] = 16'h2d1b;
initial mem[205] = 16'h2e61;
initial mem[206] = 16'h2f80;
initial mem[207] = 16'h307e;
initial mem[208] = 16'hce9f;
initial mem[209] = 16'hcf82;
initial mem[210] = 16'hd080;
initial mem[211] = 16'hd19f;
initial mem[212] = 16'hd2e5;
initial mem[213] = 16'hd459;
initial mem[214] = 16'hd606;
initial mem[215] = 16'hd7f6;
initial mem[216] = 16'hda39;
initial mem[217] = 16'hdce0;
initial mem[218] = 16'he001;
initial mem[219] = 16'he3b2;
initial mem[220] = 16'he80c;
initial mem[221] = 16'hed1d;
initial mem[222] = 16'hf2e5;
initial mem[223] = 16'hf946;
initial mem[224] = 16'h0;
initial mem[225] = 16'h5c7;
initial mem[226] = 16'hb56;
initial mem[227] = 16'h107f;
initial mem[228] = 16'h1526;
initial mem[229] = 16'h1945;
initial mem[230] = 16'h1cdf;
initial mem[231] = 16'h1fff;
initial mem[232] = 16'h22b6;
initial mem[233] = 16'h2510;
initial mem[234] = 16'h271d;
initial mem[235] = 16'h28e8;
initial mem[236] = 16'h2a7b;
initial mem[237] = 16'h2bdf;
initial mem[238] = 16'h2d1b;
initial mem[239] = 16'h2e35;
initial mem[240] = 16'hd0ce;
initial mem[241] = 16'hd1cb;
initial mem[242] = 16'hd2e5;
initial mem[243] = 16'hd421;
initial mem[244] = 16'hd585;
initial mem[245] = 16'hd718;
initial mem[246] = 16'hd8e3;
initial mem[247] = 16'hdaf0;
initial mem[248] = 16'hdd4a;
initial mem[249] = 16'he001;
initial mem[250] = 16'he321;
initial mem[251] = 16'he6bb;
initial mem[252] = 16'heada;
initial mem[253] = 16'hef81;
initial mem[254] = 16'hf4aa;
initial mem[255] = 16'hfa39;
initial mem[256] = 16'h0;
initial mem[257] = 16'h511;
initial mem[258] = 16'h9fb;
initial mem[259] = 16'he9d;
initial mem[260] = 16'h12e3;
initial mem[261] = 16'h16c2;
initial mem[262] = 16'h1a37;
initial mem[263] = 16'h1d49;
initial mem[264] = 16'h1fff;
initial mem[265] = 16'h2264;
initial mem[266] = 16'h2481;
initial mem[267] = 16'h2661;
initial mem[268] = 16'h280a;
initial mem[269] = 16'h2985;
initial mem[270] = 16'h2ad8;
initial mem[271] = 16'h2c09;
initial mem[272] = 16'hd2e5;
initial mem[273] = 16'hd3f7;
initial mem[274] = 16'hd528;
initial mem[275] = 16'hd67b;
initial mem[276] = 16'hd7f6;
initial mem[277] = 16'hd99f;
initial mem[278] = 16'hdb7f;
initial mem[279] = 16'hdd9c;
initial mem[280] = 16'he001;
initial mem[281] = 16'he2b7;
initial mem[282] = 16'he5c9;
initial mem[283] = 16'he93e;
initial mem[284] = 16'hed1d;
initial mem[285] = 16'hf163;
initial mem[286] = 16'hf605;
initial mem[287] = 16'hfaef;
initial mem[288] = 16'h0;
initial mem[289] = 16'h482;
initial mem[290] = 16'h8e8;
initial mem[291] = 16'hd1b;
initial mem[292] = 16'h110a;
initial mem[293] = 16'h14a9;
initial mem[294] = 16'h17f4;
initial mem[295] = 16'h1aee;
initial mem[296] = 16'h1d9a;
initial mem[297] = 16'h1fff;
initial mem[298] = 16'h2224;
initial mem[299] = 16'h240f;
initial mem[300] = 16'h25c7;
initial mem[301] = 16'h2753;
initial mem[302] = 16'h28b8;
initial mem[303] = 16'h29fa;
initial mem[304] = 16'hd4e1;
initial mem[305] = 16'hd606;
initial mem[306] = 16'hd748;
initial mem[307] = 16'hd8ad;
initial mem[308] = 16'hda39;
initial mem[309] = 16'hdbf1;
initial mem[310] = 16'hdddc;
initial mem[311] = 16'he001;
initial mem[312] = 16'he266;
initial mem[313] = 16'he512;
initial mem[314] = 16'he80c;
initial mem[315] = 16'heb57;
initial mem[316] = 16'heef6;
initial mem[317] = 16'hf2e5;
initial mem[318] = 16'hf718;
initial mem[319] = 16'hfb7e;
initial mem[320] = 16'h0;
initial mem[321] = 16'h40f;
initial mem[322] = 16'h80a;
initial mem[323] = 16'hbdf;
initial mem[324] = 16'hf80;
initial mem[325] = 16'h12e3;
initial mem[326] = 16'h1604;
initial mem[327] = 16'h18e1;
initial mem[328] = 16'h1b7d;
initial mem[329] = 16'h1ddb;
initial mem[330] = 16'h1fff;
initial mem[331] = 16'h21f0;
initial mem[332] = 16'h23b1;
initial mem[333] = 16'h2548;
initial mem[334] = 16'h26ba;
initial mem[335] = 16'h280a;
initial mem[336] = 16'hd6c3;
initial mem[337] = 16'hd7f6;
initial mem[338] = 16'hd946;
initial mem[339] = 16'hdab8;
initial mem[340] = 16'hdc4f;
initial mem[341] = 16'hde10;
initial mem[342] = 16'he001;
initial mem[343] = 16'he225;
initial mem[344] = 16'he483;
initial mem[345] = 16'he71f;
initial mem[346] = 16'he9fc;
initial mem[347] = 16'hed1d;
initial mem[348] = 16'hf080;
initial mem[349] = 16'hf421;
initial mem[350] = 16'hf7f6;
initial mem[351] = 16'hfbf1;
initial mem[352] = 16'h0;
initial mem[353] = 16'h3b1;
initial mem[354] = 16'h753;
initial mem[355] = 16'had9;
initial mem[356] = 16'he35;
initial mem[357] = 16'h1161;
initial mem[358] = 16'h1458;
initial mem[359] = 16'h1717;
initial mem[360] = 16'h199e;
initial mem[361] = 16'h1bf0;
initial mem[362] = 16'h1e0f;
initial mem[363] = 16'h1fff;
initial mem[364] = 16'h21c4;
initial mem[365] = 16'h2362;
initial mem[366] = 16'h24dd;
initial mem[367] = 16'h2637;
initial mem[368] = 16'hd88b;
initial mem[369] = 16'hd9c9;
initial mem[370] = 16'hdb23;
initial mem[371] = 16'hdc9e;
initial mem[372] = 16'hde3c;
initial mem[373] = 16'he001;
initial mem[374] = 16'he1f1;
initial mem[375] = 16'he410;
initial mem[376] = 16'he662;
initial mem[377] = 16'he8e9;
initial mem[378] = 16'heba8;
initial mem[379] = 16'hee9f;
initial mem[380] = 16'hf1cb;
initial mem[381] = 16'hf527;
initial mem[382] = 16'hf8ad;
initial mem[383] = 16'hfc4f;
initial mem[384] = 16'h0;
initial mem[385] = 16'h363;
initial mem[386] = 16'h6ba;
initial mem[387] = 16'h9fb;
initial mem[388] = 16'hd1b;
initial mem[389] = 16'h1015;
initial mem[390] = 16'h12e3;
initial mem[391] = 16'h1583;
initial mem[392] = 16'h17f4;
initial mem[393] = 16'h1a37;
initial mem[394] = 16'h1c4e;
initial mem[395] = 16'h1e3a;
initial mem[396] = 16'h1fff;
initial mem[397] = 16'h21a0;
initial mem[398] = 16'h2320;
initial mem[399] = 16'h2481;
initial mem[400] = 16'hda39;
initial mem[401] = 16'hdb7f;
initial mem[402] = 16'hdce0;
initial mem[403] = 16'hde60;
initial mem[404] = 16'he001;
initial mem[405] = 16'he1c6;
initial mem[406] = 16'he3b2;
initial mem[407] = 16'he5c9;
initial mem[408] = 16'he80c;
initial mem[409] = 16'hea7d;
initial mem[410] = 16'hed1d;
initial mem[411] = 16'hefeb;
initial mem[412] = 16'hf2e5;
initial mem[413] = 16'hf605;
initial mem[414] = 16'hf946;
initial mem[415] = 16'hfc9d;
initial mem[416] = 16'h0;
initial mem[417] = 16'h320;
initial mem[418] = 16'h638;
initial mem[419] = 16'h93d;
initial mem[420] = 16'hc29;
initial mem[421] = 16'hef5;
initial mem[422] = 16'h119e;
initial mem[423] = 16'h141f;
initial mem[424] = 16'h1679;
initial mem[425] = 16'h18ab;
initial mem[426] = 16'h1ab6;
initial mem[427] = 16'h1c9c;
initial mem[428] = 16'h1e5e;
initial mem[429] = 16'h1fff;
initial mem[430] = 16'h2181;
initial mem[431] = 16'h22e7;
initial mem[432] = 16'hdbce;
initial mem[433] = 16'hdd19;
initial mem[434] = 16'hde7f;
initial mem[435] = 16'he001;
initial mem[436] = 16'he1a2;
initial mem[437] = 16'he364;
initial mem[438] = 16'he54a;
initial mem[439] = 16'he755;
initial mem[440] = 16'he987;
initial mem[441] = 16'hebe1;
initial mem[442] = 16'hee62;
initial mem[443] = 16'hf10b;
initial mem[444] = 16'hf3d7;
initial mem[445] = 16'hf6c3;
initial mem[446] = 16'hf9c8;
initial mem[447] = 16'hfce0;
initial mem[448] = 16'h0;
initial mem[449] = 16'h2e7;
initial mem[450] = 16'h5c7;
initial mem[451] = 16'h899;
initial mem[452] = 16'hb56;
initial mem[453] = 16'hdf9;
initial mem[454] = 16'h107f;
initial mem[455] = 16'h12e3;
initial mem[456] = 16'h1526;
initial mem[457] = 16'h1747;
initial mem[458] = 16'h1945;
initial mem[459] = 16'h1b22;
initial mem[460] = 16'h1cdf;
initial mem[461] = 16'h1e7d;
initial mem[462] = 16'h1fff;
initial mem[463] = 16'h2167;
initial mem[464] = 16'hdd4a;
initial mem[465] = 16'hde99;
initial mem[466] = 16'he001;
initial mem[467] = 16'he183;
initial mem[468] = 16'he321;
initial mem[469] = 16'he4de;
initial mem[470] = 16'he6bb;
initial mem[471] = 16'he8b9;
initial mem[472] = 16'heada;
initial mem[473] = 16'hed1d;
initial mem[474] = 16'hef81;
initial mem[475] = 16'hf207;
initial mem[476] = 16'hf4aa;
initial mem[477] = 16'hf767;
initial mem[478] = 16'hfa39;
initial mem[479] = 16'hfd19;
initial mem[480] = 16'h0;
initial mem[481] = 16'h2b6;
initial mem[482] = 16'h566;
initial mem[483] = 16'h80a;
initial mem[484] = 16'ha9e;
initial mem[485] = 16'hd1b;
initial mem[486] = 16'hf80;
initial mem[487] = 16'h11ca;
initial mem[488] = 16'h13f6;
initial mem[489] = 16'h1604;
initial mem[490] = 16'h17f4;
initial mem[491] = 16'h19c7;
initial mem[492] = 16'h1b7d;
initial mem[493] = 16'h1d18;
initial mem[494] = 16'h1e98;
initial mem[495] = 16'h1fff;
initial mem[496] = 16'hdeb0;
initial mem[497] = 16'he001;
initial mem[498] = 16'he168;
initial mem[499] = 16'he2e8;
initial mem[500] = 16'he483;
initial mem[501] = 16'he639;
initial mem[502] = 16'he80c;
initial mem[503] = 16'he9fc;
initial mem[504] = 16'hec0a;
initial mem[505] = 16'hee36;
initial mem[506] = 16'hf080;
initial mem[507] = 16'hf2e5;
initial mem[508] = 16'hf562;
initial mem[509] = 16'hf7f6;
initial mem[510] = 16'hfa9a;
initial mem[511] = 16'hfd4a;
initial mem[512] = 16'h7fff;
initial mem[513] = 16'h7d73;
initial mem[514] = 16'h7aed;
initial mem[515] = 16'h7871;
initial mem[516] = 16'h7603;
initial mem[517] = 16'h73a7;
initial mem[518] = 16'h7161;
initial mem[519] = 16'h6f31;
initial mem[520] = 16'h6d1b;
initial mem[521] = 16'h6b1e;
initial mem[522] = 16'h693c;
initial mem[523] = 16'h6775;
initial mem[524] = 16'h65c7;
initial mem[525] = 16'h6432;
initial mem[526] = 16'h62b5;
initial mem[527] = 16'h614f;
initial mem[528] = 16'ha001;
initial mem[529] = 16'h9eb1;
initial mem[530] = 16'h9d4b;
initial mem[531] = 16'h9bce;
initial mem[532] = 16'h9a39;
initial mem[533] = 16'h988b;
initial mem[534] = 16'h96c4;
initial mem[535] = 16'h94e2;
initial mem[536] = 16'h92e5;
initial mem[537] = 16'h90cf;
initial mem[538] = 16'h8e9f;
initial mem[539] = 16'h8c59;
initial mem[540] = 16'h89fd;
initial mem[541] = 16'h878f;
initial mem[542] = 16'h8513;
initial mem[543] = 16'h828d;
initial mem[544] = 16'h7fff;
initial mem[545] = 16'h7d48;
initial mem[546] = 16'h7a98;
initial mem[547] = 16'h77f4;
initial mem[548] = 16'h7560;
initial mem[549] = 16'h72e3;
initial mem[550] = 16'h707e;
initial mem[551] = 16'h6e34;
initial mem[552] = 16'h6c08;
initial mem[553] = 16'h69fa;
initial mem[554] = 16'h680a;
initial mem[555] = 16'h6637;
initial mem[556] = 16'h6481;
initial mem[557] = 16'h62e6;
initial mem[558] = 16'h6166;
initial mem[559] = 16'h5fff;
initial mem[560] = 16'ha152;
initial mem[561] = 16'ha001;
initial mem[562] = 16'h9e9a;
initial mem[563] = 16'h9d1a;
initial mem[564] = 16'h9b7f;
initial mem[565] = 16'h99c9;
initial mem[566] = 16'h97f6;
initial mem[567] = 16'h9606;
initial mem[568] = 16'h93f8;
initial mem[569] = 16'h91cc;
initial mem[570] = 16'h8f82;
initial mem[571] = 16'h8d1d;
initial mem[572] = 16'h8aa0;
initial mem[573] = 16'h880c;
initial mem[574] = 16'h8568;
initial mem[575] = 16'h82b8;
initial mem[576] = 16'h7fff;
initial mem[577] = 16'h7d17;
initial mem[578] = 16'h7a37;
initial mem[579] = 16'h7765;
initial mem[580] = 16'h74a8;
initial mem[581] = 16'h7205;
initial mem[582] = 16'h6f7f;
initial mem[583] = 16'h6d1b;
initial mem[584] = 16'h6ad8;
initial mem[585] = 16'h68b7;
initial mem[586] = 16'h66b9;
initial mem[587] = 16'h64dc;
initial mem[588] = 16'h631f;
initial mem[589] = 16'h6181;
initial mem[590] = 16'h5fff;
initial mem[591] = 16'h5e97;
initial mem[592] = 16'ha2b8;
initial mem[593] = 16'ha169;
initial mem[594] = 16'ha001;
initial mem[595] = 16'h9e7f;
initial mem[596] = 16'h9ce1;
initial mem[597] = 16'h9b24;
initial mem[598] = 16'h9947;
initial mem[599] = 16'h9749;
initial mem[600] = 16'h9528;
initial mem[601] = 16'h92e5;
initial mem[602] = 16'h9081;
initial mem[603] = 16'h8dfb;
initial mem[604] = 16'h8b58;
initial mem[605] = 16'h889b;
initial mem[606] = 16'h85c9;
initial mem[607] = 16'h82e9;
initial mem[608] = 16'h7fff;
initial mem[609] = 16'h7cde;
initial mem[610] = 16'h79c6;
initial mem[611] = 16'h76c1;
initial mem[612] = 16'h73d5;
initial mem[613] = 16'h7109;
initial mem[614] = 16'h6e60;
initial mem[615] = 16'h6bdf;
initial mem[616] = 16'h6985;
initial mem[617] = 16'h6753;
initial mem[618] = 16'h6548;
initial mem[619] = 16'h6362;
initial mem[620] = 16'h61a0;
initial mem[621] = 16'h5fff;
initial mem[622] = 16'h5e7d;
initial mem[623] = 16'h5d17;
initial mem[624] = 16'ha434;
initial mem[625] = 16'ha2e9;
initial mem[626] = 16'ha183;
initial mem[627] = 16'ha001;
initial mem[628] = 16'h9e60;
initial mem[629] = 16'h9c9e;
initial mem[630] = 16'h9ab8;
initial mem[631] = 16'h98ad;
initial mem[632] = 16'h967b;
initial mem[633] = 16'h9421;
initial mem[634] = 16'h91a0;
initial mem[635] = 16'h8ef7;
initial mem[636] = 16'h8c2b;
initial mem[637] = 16'h893f;
initial mem[638] = 16'h863a;
initial mem[639] = 16'h8322;
initial mem[640] = 16'h7fff;
initial mem[641] = 16'h7c9b;
initial mem[642] = 16'h7944;
initial mem[643] = 16'h7603;
initial mem[644] = 16'h72e3;
initial mem[645] = 16'h6fe9;
initial mem[646] = 16'h6d1b;
initial mem[647] = 16'h6a7b;
initial mem[648] = 16'h680a;
initial mem[649] = 16'h65c7;
initial mem[650] = 16'h63b0;
initial mem[651] = 16'h61c4;
initial mem[652] = 16'h5fff;
initial mem[653] = 16'h5e5e;
initial mem[654] = 16'h5cde;
initial mem[655] = 16'h5b7d;
initial mem[656] = 16'ha5c9;
initial mem[657] = 16'ha483;
initial mem[658] = 16'ha322;
initial mem[659] = 16'ha1a2;
initial mem[660] = 16'ha001;
initial mem[661] = 16'h9e3c;
initial mem[662] = 16'h9c50;
initial mem[663] = 16'h9a39;
initial mem[664] = 16'h97f6;
initial mem[665] = 16'h9585;
initial mem[666] = 16'h92e5;
initial mem[667] = 16'h9017;
initial mem[668] = 16'h8d1d;
initial mem[669] = 16'h89fd;
initial mem[670] = 16'h86bc;
initial mem[671] = 16'h8365;
initial mem[672] = 16'h7fff;
initial mem[673] = 16'h7c4d;
initial mem[674] = 16'h78ab;
initial mem[675] = 16'h7525;
initial mem[676] = 16'h71c9;
initial mem[677] = 16'h6e9d;
initial mem[678] = 16'h6ba6;
initial mem[679] = 16'h68e7;
initial mem[680] = 16'h6660;
initial mem[681] = 16'h640e;
initial mem[682] = 16'h61ef;
initial mem[683] = 16'h5fff;
initial mem[684] = 16'h5e3a;
initial mem[685] = 16'h5c9c;
initial mem[686] = 16'h5b21;
initial mem[687] = 16'h59c7;
initial mem[688] = 16'ha777;
initial mem[689] = 16'ha639;
initial mem[690] = 16'ha4df;
initial mem[691] = 16'ha364;
initial mem[692] = 16'ha1c6;
initial mem[693] = 16'ha001;
initial mem[694] = 16'h9e11;
initial mem[695] = 16'h9bf2;
initial mem[696] = 16'h99a0;
initial mem[697] = 16'h9719;
initial mem[698] = 16'h945a;
initial mem[699] = 16'h9163;
initial mem[700] = 16'h8e37;
initial mem[701] = 16'h8adb;
initial mem[702] = 16'h8755;
initial mem[703] = 16'h83b3;
initial mem[704] = 16'h7fff;
initial mem[705] = 16'h7bef;
initial mem[706] = 16'h77f4;
initial mem[707] = 16'h741f;
initial mem[708] = 16'h707e;
initial mem[709] = 16'h6d1b;
initial mem[710] = 16'h69fa;
initial mem[711] = 16'h671d;
initial mem[712] = 16'h6481;
initial mem[713] = 16'h6223;
initial mem[714] = 16'h5fff;
initial mem[715] = 16'h5e0e;
initial mem[716] = 16'h5c4d;
initial mem[717] = 16'h5ab6;
initial mem[718] = 16'h5944;
initial mem[719] = 16'h57f4;
initial mem[720] = 16'ha93f;
initial mem[721] = 16'ha80c;
initial mem[722] = 16'ha6bc;
initial mem[723] = 16'ha54a;
initial mem[724] = 16'ha3b3;
initial mem[725] = 16'ha1f2;
initial mem[726] = 16'ha001;
initial mem[727] = 16'h9ddd;
initial mem[728] = 16'h9b7f;
initial mem[729] = 16'h98e3;
initial mem[730] = 16'h9606;
initial mem[731] = 16'h92e5;
initial mem[732] = 16'h8f82;
initial mem[733] = 16'h8be1;
initial mem[734] = 16'h880c;
initial mem[735] = 16'h8411;
initial mem[736] = 16'h7fff;
initial mem[737] = 16'h7b7c;
initial mem[738] = 16'h7716;
initial mem[739] = 16'h72e3;
initial mem[740] = 16'h6ef4;
initial mem[741] = 16'h6b55;
initial mem[742] = 16'h680a;
initial mem[743] = 16'h6510;
initial mem[744] = 16'h6264;
initial mem[745] = 16'h5fff;
initial mem[746] = 16'h5dda;
initial mem[747] = 16'h5bef;
initial mem[748] = 16'h5a37;
initial mem[749] = 16'h58ab;
initial mem[750] = 16'h5746;
initial mem[751] = 16'h5604;
initial mem[752] = 16'hab21;
initial mem[753] = 16'ha9fc;
initial mem[754] = 16'ha8ba;
initial mem[755] = 16'ha755;
initial mem[756] = 16'ha5c9;
initial mem[757] = 16'ha411;
initial mem[758] = 16'ha226;
initial mem[759] = 16'ha001;
initial mem[760] = 16'h9d9c;
initial mem[761] = 16'h9af0;
initial mem[762] = 16'h97f6;
initial mem[763] = 16'h94ab;
initial mem[764] = 16'h910c;
initial mem[765] = 16'h8d1d;
initial mem[766] = 16'h88ea;
initial mem[767] = 16'h8484;
initial mem[768] = 16'h7fff;
initial mem[769] = 16'h7aed;
initial mem[770] = 16'h7603;
initial mem[771] = 16'h7161;
initial mem[772] = 16'h6d1b;
initial mem[773] = 16'h693c;
initial mem[774] = 16'h65c7;
initial mem[775] = 16'h62b5;
initial mem[776] = 16'h5fff;
initial mem[777] = 16'h5d9a;
initial mem[778] = 16'h5b7d;
initial mem[779] = 16'h599d;
initial mem[780] = 16'h57f4;
initial mem[781] = 16'h5679;
initial mem[782] = 16'h5526;
initial mem[783] = 16'h53f5;
initial mem[784] = 16'had1d;
initial mem[785] = 16'hac0b;
initial mem[786] = 16'haada;
initial mem[787] = 16'ha987;
initial mem[788] = 16'ha80c;
initial mem[789] = 16'ha663;
initial mem[790] = 16'ha483;
initial mem[791] = 16'ha266;
initial mem[792] = 16'ha001;
initial mem[793] = 16'h9d4b;
initial mem[794] = 16'h9a39;
initial mem[795] = 16'h96c4;
initial mem[796] = 16'h92e5;
initial mem[797] = 16'h8e9f;
initial mem[798] = 16'h89fd;
initial mem[799] = 16'h8513;
initial mem[800] = 16'h7fff;
initial mem[801] = 16'h7a37;
initial mem[802] = 16'h74a8;
initial mem[803] = 16'h6f7f;
initial mem[804] = 16'h6ad8;
initial mem[805] = 16'h66b9;
initial mem[806] = 16'h631f;
initial mem[807] = 16'h5fff;
initial mem[808] = 16'h5d48;
initial mem[809] = 16'h5aee;
initial mem[810] = 16'h58e1;
initial mem[811] = 16'h5716;
initial mem[812] = 16'h5583;
initial mem[813] = 16'h541f;
initial mem[814] = 16'h52e3;
initial mem[815] = 16'h51c9;
initial mem[816] = 16'haf34;
initial mem[817] = 16'hae37;
initial mem[818] = 16'had1d;
initial mem[819] = 16'habe1;
initial mem[820] = 16'haa7d;
initial mem[821] = 16'ha8ea;
initial mem[822] = 16'ha71f;
initial mem[823] = 16'ha512;
initial mem[824] = 16'ha2b8;
initial mem[825] = 16'ha001;
initial mem[826] = 16'h9ce1;
initial mem[827] = 16'h9947;
initial mem[828] = 16'h9528;
initial mem[829] = 16'h9081;
initial mem[830] = 16'h8b58;
initial mem[831] = 16'h85c9;
initial mem[832] = 16'h7fff;
initial mem[833] = 16'h7944;
initial mem[834] = 16'h72e3;
initial mem[835] = 16'h6d1b;
initial mem[836] = 16'h680a;
initial mem[837] = 16'h63b0;
initial mem[838] = 16'h5fff;
initial mem[839] = 16'h5cde;
initial mem[840] = 16'h5a37;
initial mem[841] = 16'h57f4;
initial mem[842] = 16'h5604;
initial mem[843] = 16'h5457;
initial mem[844] = 16'h52e3;
initial mem[845] = 16'h519d;
initial mem[846] = 16'h507e;
initial mem[847] = 16'h4f80;
initial mem[848] = 16'hb163;
initial mem[849] = 16'hb080;
initial mem[850] = 16'haf82;
initial mem[851] = 16'hae63;
initial mem[852] = 16'had1d;
initial mem[853] = 16'haba9;
initial mem[854] = 16'ha9fc;
initial mem[855] = 16'ha80c;
initial mem[856] = 16'ha5c9;
initial mem[857] = 16'ha322;
initial mem[858] = 16'ha001;
initial mem[859] = 16'h9c50;
initial mem[860] = 16'h97f6;
initial mem[861] = 16'h92e5;
initial mem[862] = 16'h8d1d;
initial mem[863] = 16'h86bc;
initial mem[864] = 16'h7fff;
initial mem[865] = 16'h77f4;
initial mem[866] = 16'h707e;
initial mem[867] = 16'h69fa;
initial mem[868] = 16'h6481;
initial mem[869] = 16'h5fff;
initial mem[870] = 16'h5c4d;
initial mem[871] = 16'h5944;
initial mem[872] = 16'h56c1;
initial mem[873] = 16'h54a8;
initial mem[874] = 16'h52e3;
initial mem[875] = 16'h5161;
initial mem[876] = 16'h5015;
initial mem[877] = 16'h4ef5;
initial mem[878] = 16'h4df9;
initial mem[879] = 16'h4d1b;
initial mem[880] = 16'hb3aa;
initial mem[881] = 16'hb2e5;
initial mem[882] = 16'hb207;
initial mem[883] = 16'hb10b;
initial mem[884] = 16'hafeb;
initial mem[885] = 16'hae9f;
initial mem[886] = 16'had1d;
initial mem[887] = 16'hab58;
initial mem[888] = 16'ha93f;
initial mem[889] = 16'ha6bc;
initial mem[890] = 16'ha3b3;
initial mem[891] = 16'ha001;
initial mem[892] = 16'h9b7f;
initial mem[893] = 16'h9606;
initial mem[894] = 16'h8f82;
initial mem[895] = 16'h880c;
initial mem[896] = 16'h7fff;
initial mem[897] = 16'h7603;
initial mem[898] = 16'h6d1b;
initial mem[899] = 16'h65c7;
initial mem[900] = 16'h5fff;
initial mem[901] = 16'h5b7d;
initial mem[902] = 16'h57f4;
initial mem[903] = 16'h5526;
initial mem[904] = 16'h52e3;
initial mem[905] = 16'h5109;
initial mem[906] = 16'h4f80;
initial mem[907] = 16'h4e35;
initial mem[908] = 16'h4d1b;
initial mem[909] = 16'h4c28;
initial mem[910] = 16'h4b56;
initial mem[911] = 16'h4a9d;
initial mem[912] = 16'hb606;
initial mem[913] = 16'hb563;
initial mem[914] = 16'hb4aa;
initial mem[915] = 16'hb3d8;
initial mem[916] = 16'hb2e5;
initial mem[917] = 16'hb1cb;
initial mem[918] = 16'hb080;
initial mem[919] = 16'haef7;
initial mem[920] = 16'had1d;
initial mem[921] = 16'haada;
initial mem[922] = 16'ha80c;
initial mem[923] = 16'ha483;
initial mem[924] = 16'ha001;
initial mem[925] = 16'h9a39;
initial mem[926] = 16'h92e5;
initial mem[927] = 16'h89fd;
initial mem[928] = 16'h7fff;
initial mem[929] = 16'h72e3;
initial mem[930] = 16'h680a;
initial mem[931] = 16'h5fff;
initial mem[932] = 16'h5a37;
initial mem[933] = 16'h5604;
initial mem[934] = 16'h52e3;
initial mem[935] = 16'h507e;
initial mem[936] = 16'h4e9d;
initial mem[937] = 16'h4d1b;
initial mem[938] = 16'h4bdf;
initial mem[939] = 16'h4ad8;
initial mem[940] = 16'h49fa;
initial mem[941] = 16'h493d;
initial mem[942] = 16'h4899;
initial mem[943] = 16'h480a;
initial mem[944] = 16'hb874;
initial mem[945] = 16'hb7f6;
initial mem[946] = 16'hb767;
initial mem[947] = 16'hb6c3;
initial mem[948] = 16'hb606;
initial mem[949] = 16'hb528;
initial mem[950] = 16'hb421;
initial mem[951] = 16'hb2e5;
initial mem[952] = 16'hb163;
initial mem[953] = 16'haf82;
initial mem[954] = 16'had1d;
initial mem[955] = 16'ha9fc;
initial mem[956] = 16'ha5c9;
initial mem[957] = 16'ha001;
initial mem[958] = 16'h97f6;
initial mem[959] = 16'h8d1d;
initial mem[960] = 16'h7fff;
initial mem[961] = 16'h6d1b;
initial mem[962] = 16'h5fff;
initial mem[963] = 16'h57f4;
initial mem[964] = 16'h52e3;
initial mem[965] = 16'h4f80;
initial mem[966] = 16'h4d1b;
initial mem[967] = 16'h4b56;
initial mem[968] = 16'h49fa;
initial mem[969] = 16'h48e8;
initial mem[970] = 16'h480a;
initial mem[971] = 16'h4753;
initial mem[972] = 16'h46ba;
initial mem[973] = 16'h4637;
initial mem[974] = 16'h45c7;
initial mem[975] = 16'h4566;
initial mem[976] = 16'hbaf0;
initial mem[977] = 16'hba9a;
initial mem[978] = 16'hba39;
initial mem[979] = 16'hb9c9;
initial mem[980] = 16'hb946;
initial mem[981] = 16'hb8ad;
initial mem[982] = 16'hb7f6;
initial mem[983] = 16'hb718;
initial mem[984] = 16'hb606;
initial mem[985] = 16'hb4aa;
initial mem[986] = 16'hb2e5;
initial mem[987] = 16'hb080;
initial mem[988] = 16'had1d;
initial mem[989] = 16'ha80c;
initial mem[990] = 16'ha001;
initial mem[991] = 16'h92e5;
initial mem[992] = 16'h7fff;
initial mem[993] = 16'h5fff;
initial mem[994] = 16'h52e3;
initial mem[995] = 16'h4d1b;
initial mem[996] = 16'h49fa;
initial mem[997] = 16'h480a;
initial mem[998] = 16'h46ba;
initial mem[999] = 16'h45c7;
initial mem[1000] = 16'h4510;
initial mem[1001] = 16'h4481;
initial mem[1002] = 16'h440f;
initial mem[1003] = 16'h43b1;
initial mem[1004] = 16'h4362;
initial mem[1005] = 16'h4320;
initial mem[1006] = 16'h42e7;
initial mem[1007] = 16'h42b5;
initial mem[1008] = 16'hbd76;
initial mem[1009] = 16'hbd4b;
initial mem[1010] = 16'hbd19;
initial mem[1011] = 16'hbce0;
initial mem[1012] = 16'hbc9e;
initial mem[1013] = 16'hbc4f;
initial mem[1014] = 16'hbbf1;
initial mem[1015] = 16'hbb7f;
initial mem[1016] = 16'hbaf0;
initial mem[1017] = 16'hba39;
initial mem[1018] = 16'hb946;
initial mem[1019] = 16'hb7f6;
initial mem[1020] = 16'hb606;
initial mem[1021] = 16'hb2e5;
initial mem[1022] = 16'had1d;
initial mem[1023] = 16'ha001;
always @(posedge clk) begin
	data <= mem[addr];
end
endmodule
