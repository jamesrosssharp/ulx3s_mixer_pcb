module argTable(input clk, input [9:0] addr, output reg [15:0] data);
reg [15:0] mem [0:1023];
initial mem[0] = 16'h0;
initial mem[1] = 16'h7fff;
initial mem[2] = 16'h7fff;
initial mem[3] = 16'h7fff;
initial mem[4] = 16'h7fff;
initial mem[5] = 16'h7fff;
initial mem[6] = 16'h7fff;
initial mem[7] = 16'h7fff;
initial mem[8] = 16'h7fff;
initial mem[9] = 16'h7fff;
initial mem[10] = 16'h7fff;
initial mem[11] = 16'h7fff;
initial mem[12] = 16'h7fff;
initial mem[13] = 16'h7fff;
initial mem[14] = 16'h7fff;
initial mem[15] = 16'h7fff;
initial mem[16] = 16'h8001;
initial mem[17] = 16'h8001;
initial mem[18] = 16'h8001;
initial mem[19] = 16'h8001;
initial mem[20] = 16'h8001;
initial mem[21] = 16'h8001;
initial mem[22] = 16'h8001;
initial mem[23] = 16'h8001;
initial mem[24] = 16'h8001;
initial mem[25] = 16'h8001;
initial mem[26] = 16'h8001;
initial mem[27] = 16'h8001;
initial mem[28] = 16'h8001;
initial mem[29] = 16'h8001;
initial mem[30] = 16'h8001;
initial mem[31] = 16'h8001;
initial mem[32] = 16'h0;
initial mem[33] = 16'h3fff;
initial mem[34] = 16'h5a37;
initial mem[35] = 16'h65c7;
initial mem[36] = 16'h6c08;
initial mem[37] = 16'h6fe9;
initial mem[38] = 16'h7289;
initial mem[39] = 16'h746f;
initial mem[40] = 16'h75dc;
initial mem[41] = 16'h76fa;
initial mem[42] = 16'h77df;
initial mem[43] = 16'h789b;
initial mem[44] = 16'h7938;
initial mem[45] = 16'h79bd;
initial mem[46] = 16'h7a2f;
initial mem[47] = 16'h7a92;
initial mem[48] = 16'h8518;
initial mem[49] = 16'h856e;
initial mem[50] = 16'h85d1;
initial mem[51] = 16'h8643;
initial mem[52] = 16'h86c8;
initial mem[53] = 16'h8765;
initial mem[54] = 16'h8821;
initial mem[55] = 16'h8906;
initial mem[56] = 16'h8a24;
initial mem[57] = 16'h8b91;
initial mem[58] = 16'h8d77;
initial mem[59] = 16'h9017;
initial mem[60] = 16'h93f8;
initial mem[61] = 16'h9a39;
initial mem[62] = 16'ha5c9;
initial mem[63] = 16'hc001;
initial mem[64] = 16'h0;
initial mem[65] = 16'h25c7;
initial mem[66] = 16'h3fff;
initial mem[67] = 16'h5015;
initial mem[68] = 16'h5a37;
initial mem[69] = 16'h60fd;
initial mem[70] = 16'h65c7;
initial mem[71] = 16'h6951;
initial mem[72] = 16'h6c08;
initial mem[73] = 16'h6e2d;
initial mem[74] = 16'h6fe9;
initial mem[75] = 16'h7157;
initial mem[76] = 16'h7289;
initial mem[77] = 16'h738e;
initial mem[78] = 16'h746f;
initial mem[79] = 16'h7531;
initial mem[80] = 16'h8a24;
initial mem[81] = 16'h8acf;
initial mem[82] = 16'h8b91;
initial mem[83] = 16'h8c72;
initial mem[84] = 16'h8d77;
initial mem[85] = 16'h8ea9;
initial mem[86] = 16'h9017;
initial mem[87] = 16'h91d3;
initial mem[88] = 16'h93f8;
initial mem[89] = 16'h96af;
initial mem[90] = 16'h9a39;
initial mem[91] = 16'h9f03;
initial mem[92] = 16'ha5c9;
initial mem[93] = 16'hafeb;
initial mem[94] = 16'hc001;
initial mem[95] = 16'hda39;
initial mem[96] = 16'h0;
initial mem[97] = 16'h1a37;
initial mem[98] = 16'h2fe9;
initial mem[99] = 16'h3fff;
initial mem[100] = 16'h4b8f;
initial mem[101] = 16'h53f5;
initial mem[102] = 16'h5a37;
initial mem[103] = 16'h5f00;
initial mem[104] = 16'h62c3;
initial mem[105] = 16'h65c7;
initial mem[106] = 16'h683f;
initial mem[107] = 16'h6a4c;
initial mem[108] = 16'h6c08;
initial mem[109] = 16'h6d83;
initial mem[110] = 16'h6ecb;
initial mem[111] = 16'h6fe9;
initial mem[112] = 16'h8f1c;
initial mem[113] = 16'h9017;
initial mem[114] = 16'h9135;
initial mem[115] = 16'h927d;
initial mem[116] = 16'h93f8;
initial mem[117] = 16'h95b4;
initial mem[118] = 16'h97c1;
initial mem[119] = 16'h9a39;
initial mem[120] = 16'h9d3d;
initial mem[121] = 16'ha100;
initial mem[122] = 16'ha5c9;
initial mem[123] = 16'hac0b;
initial mem[124] = 16'hb471;
initial mem[125] = 16'hc001;
initial mem[126] = 16'hd017;
initial mem[127] = 16'he5c9;
initial mem[128] = 16'h0;
initial mem[129] = 16'h13f6;
initial mem[130] = 16'h25c7;
initial mem[131] = 16'h346f;
initial mem[132] = 16'h3fff;
initial mem[133] = 16'h4903;
initial mem[134] = 16'h5015;
initial mem[135] = 16'h55b1;
initial mem[136] = 16'h5a37;
initial mem[137] = 16'h5dea;
initial mem[138] = 16'h60fd;
initial mem[139] = 16'h6393;
initial mem[140] = 16'h65c7;
initial mem[141] = 16'h67ac;
initial mem[142] = 16'h6951;
initial mem[143] = 16'h6ac2;
initial mem[144] = 16'h93f8;
initial mem[145] = 16'h953e;
initial mem[146] = 16'h96af;
initial mem[147] = 16'h9854;
initial mem[148] = 16'h9a39;
initial mem[149] = 16'h9c6d;
initial mem[150] = 16'h9f03;
initial mem[151] = 16'ha216;
initial mem[152] = 16'ha5c9;
initial mem[153] = 16'haa4f;
initial mem[154] = 16'hafeb;
initial mem[155] = 16'hb6fd;
initial mem[156] = 16'hc001;
initial mem[157] = 16'hcb91;
initial mem[158] = 16'hda39;
initial mem[159] = 16'hec0a;
initial mem[160] = 16'h0;
initial mem[161] = 16'h1015;
initial mem[162] = 16'h1f01;
initial mem[163] = 16'h2c09;
initial mem[164] = 16'h36fb;
initial mem[165] = 16'h3fff;
initial mem[166] = 16'h4762;
initial mem[167] = 16'h4d74;
initial mem[168] = 16'h527a;
initial mem[169] = 16'h56ac;
initial mem[170] = 16'h5a37;
initial mem[171] = 16'h5d3b;
initial mem[172] = 16'h5fd3;
initial mem[173] = 16'h6213;
initial mem[174] = 16'h640b;
initial mem[175] = 16'h65c7;
initial mem[176] = 16'h98b0;
initial mem[177] = 16'h9a39;
initial mem[178] = 16'h9bf5;
initial mem[179] = 16'h9ded;
initial mem[180] = 16'ha02d;
initial mem[181] = 16'ha2c5;
initial mem[182] = 16'ha5c9;
initial mem[183] = 16'ha954;
initial mem[184] = 16'had86;
initial mem[185] = 16'hb28c;
initial mem[186] = 16'hb89e;
initial mem[187] = 16'hc001;
initial mem[188] = 16'hc905;
initial mem[189] = 16'hd3f7;
initial mem[190] = 16'he0ff;
initial mem[191] = 16'hefeb;
initial mem[192] = 16'h0;
initial mem[193] = 16'hd75;
initial mem[194] = 16'h1a37;
initial mem[195] = 16'h25c7;
initial mem[196] = 16'h2fe9;
initial mem[197] = 16'h389c;
initial mem[198] = 16'h3fff;
initial mem[199] = 16'h4640;
initial mem[200] = 16'h4b8f;
initial mem[201] = 16'h5015;
initial mem[202] = 16'h53f5;
initial mem[203] = 16'h574e;
initial mem[204] = 16'h5a37;
initial mem[205] = 16'h5cc2;
initial mem[206] = 16'h5f00;
initial mem[207] = 16'h60fd;
initial mem[208] = 16'h9d3d;
initial mem[209] = 16'h9f03;
initial mem[210] = 16'ha100;
initial mem[211] = 16'ha33e;
initial mem[212] = 16'ha5c9;
initial mem[213] = 16'ha8b2;
initial mem[214] = 16'hac0b;
initial mem[215] = 16'hafeb;
initial mem[216] = 16'hb471;
initial mem[217] = 16'hb9c0;
initial mem[218] = 16'hc001;
initial mem[219] = 16'hc764;
initial mem[220] = 16'hd017;
initial mem[221] = 16'hda39;
initial mem[222] = 16'he5c9;
initial mem[223] = 16'hf28b;
initial mem[224] = 16'h0;
initial mem[225] = 16'hb8f;
initial mem[226] = 16'h16ad;
initial mem[227] = 16'h20fe;
initial mem[228] = 16'h2a4d;
initial mem[229] = 16'h328a;
initial mem[230] = 16'h39be;
initial mem[231] = 16'h3fff;
initial mem[232] = 16'h456c;
initial mem[233] = 16'h4a21;
initial mem[234] = 16'h4e3b;
initial mem[235] = 16'h51d0;
initial mem[236] = 16'h54f7;
initial mem[237] = 16'h57bf;
initial mem[238] = 16'h5a37;
initial mem[239] = 16'h5c6a;
initial mem[240] = 16'ha19c;
initial mem[241] = 16'ha396;
initial mem[242] = 16'ha5c9;
initial mem[243] = 16'ha841;
initial mem[244] = 16'hab09;
initial mem[245] = 16'hae30;
initial mem[246] = 16'hb1c5;
initial mem[247] = 16'hb5df;
initial mem[248] = 16'hba94;
initial mem[249] = 16'hc001;
initial mem[250] = 16'hc642;
initial mem[251] = 16'hcd76;
initial mem[252] = 16'hd5b3;
initial mem[253] = 16'hdf02;
initial mem[254] = 16'he953;
initial mem[255] = 16'hf471;
initial mem[256] = 16'h0;
initial mem[257] = 16'ha22;
initial mem[258] = 16'h13f6;
initial mem[259] = 16'h1d3b;
initial mem[260] = 16'h25c7;
initial mem[261] = 16'h2d84;
initial mem[262] = 16'h346f;
initial mem[263] = 16'h3a92;
initial mem[264] = 16'h3fff;
initial mem[265] = 16'h44c9;
initial mem[266] = 16'h4903;
initial mem[267] = 16'h4cc2;
initial mem[268] = 16'h5015;
initial mem[269] = 16'h530b;
initial mem[270] = 16'h55b1;
initial mem[271] = 16'h5812;
initial mem[272] = 16'ha5c9;
initial mem[273] = 16'ha7ee;
initial mem[274] = 16'haa4f;
initial mem[275] = 16'hacf5;
initial mem[276] = 16'hafeb;
initial mem[277] = 16'hb33e;
initial mem[278] = 16'hb6fd;
initial mem[279] = 16'hbb37;
initial mem[280] = 16'hc001;
initial mem[281] = 16'hc56e;
initial mem[282] = 16'hcb91;
initial mem[283] = 16'hd27c;
initial mem[284] = 16'hda39;
initial mem[285] = 16'he2c5;
initial mem[286] = 16'hec0a;
initial mem[287] = 16'hf5de;
initial mem[288] = 16'h0;
initial mem[289] = 16'h904;
initial mem[290] = 16'h11d1;
initial mem[291] = 16'h1a37;
initial mem[292] = 16'h2214;
initial mem[293] = 16'h2952;
initial mem[294] = 16'h2fe9;
initial mem[295] = 16'h35dd;
initial mem[296] = 16'h3b35;
initial mem[297] = 16'h3fff;
initial mem[298] = 16'h4448;
initial mem[299] = 16'h481e;
initial mem[300] = 16'h4b8f;
initial mem[301] = 16'h4ea7;
initial mem[302] = 16'h5170;
initial mem[303] = 16'h53f5;
initial mem[304] = 16'ha9c2;
initial mem[305] = 16'hac0b;
initial mem[306] = 16'hae90;
initial mem[307] = 16'hb159;
initial mem[308] = 16'hb471;
initial mem[309] = 16'hb7e2;
initial mem[310] = 16'hbbb8;
initial mem[311] = 16'hc001;
initial mem[312] = 16'hc4cb;
initial mem[313] = 16'hca23;
initial mem[314] = 16'hd017;
initial mem[315] = 16'hd6ae;
initial mem[316] = 16'hddec;
initial mem[317] = 16'he5c9;
initial mem[318] = 16'hee2f;
initial mem[319] = 16'hf6fc;
initial mem[320] = 16'h0;
initial mem[321] = 16'h81f;
initial mem[322] = 16'h1015;
initial mem[323] = 16'h17bf;
initial mem[324] = 16'h1f01;
initial mem[325] = 16'h25c7;
initial mem[326] = 16'h2c09;
initial mem[327] = 16'h31c3;
initial mem[328] = 16'h36fb;
initial mem[329] = 16'h3bb6;
initial mem[330] = 16'h3fff;
initial mem[331] = 16'h43e0;
initial mem[332] = 16'h4762;
initial mem[333] = 16'h4a91;
initial mem[334] = 16'h4d74;
initial mem[335] = 16'h5015;
initial mem[336] = 16'had86;
initial mem[337] = 16'hafeb;
initial mem[338] = 16'hb28c;
initial mem[339] = 16'hb56f;
initial mem[340] = 16'hb89e;
initial mem[341] = 16'hbc20;
initial mem[342] = 16'hc001;
initial mem[343] = 16'hc44a;
initial mem[344] = 16'hc905;
initial mem[345] = 16'hce3d;
initial mem[346] = 16'hd3f7;
initial mem[347] = 16'hda39;
initial mem[348] = 16'he0ff;
initial mem[349] = 16'he841;
initial mem[350] = 16'hefeb;
initial mem[351] = 16'hf7e1;
initial mem[352] = 16'h0;
initial mem[353] = 16'h763;
initial mem[354] = 16'hea7;
initial mem[355] = 16'h15b2;
initial mem[356] = 16'h1c6b;
initial mem[357] = 16'h22c3;
initial mem[358] = 16'h28b0;
initial mem[359] = 16'h2e2e;
initial mem[360] = 16'h333c;
initial mem[361] = 16'h37e0;
initial mem[362] = 16'h3c1e;
initial mem[363] = 16'h3fff;
initial mem[364] = 16'h4389;
initial mem[365] = 16'h46c5;
initial mem[366] = 16'h49ba;
initial mem[367] = 16'h4c6f;
initial mem[368] = 16'hb115;
initial mem[369] = 16'hb391;
initial mem[370] = 16'hb646;
initial mem[371] = 16'hb93b;
initial mem[372] = 16'hbc77;
initial mem[373] = 16'hc001;
initial mem[374] = 16'hc3e2;
initial mem[375] = 16'hc820;
initial mem[376] = 16'hccc4;
initial mem[377] = 16'hd1d2;
initial mem[378] = 16'hd750;
initial mem[379] = 16'hdd3d;
initial mem[380] = 16'he395;
initial mem[381] = 16'hea4e;
initial mem[382] = 16'hf159;
initial mem[383] = 16'hf89d;
initial mem[384] = 16'h0;
initial mem[385] = 16'h6c6;
initial mem[386] = 16'hd75;
initial mem[387] = 16'h13f6;
initial mem[388] = 16'h1a37;
initial mem[389] = 16'h202b;
initial mem[390] = 16'h25c7;
initial mem[391] = 16'h2b07;
initial mem[392] = 16'h2fe9;
initial mem[393] = 16'h346f;
initial mem[394] = 16'h389c;
initial mem[395] = 16'h3c75;
initial mem[396] = 16'h3fff;
initial mem[397] = 16'h4341;
initial mem[398] = 16'h4640;
initial mem[399] = 16'h4903;
initial mem[400] = 16'hb471;
initial mem[401] = 16'hb6fd;
initial mem[402] = 16'hb9c0;
initial mem[403] = 16'hbcbf;
initial mem[404] = 16'hc001;
initial mem[405] = 16'hc38b;
initial mem[406] = 16'hc764;
initial mem[407] = 16'hcb91;
initial mem[408] = 16'hd017;
initial mem[409] = 16'hd4f9;
initial mem[410] = 16'hda39;
initial mem[411] = 16'hdfd5;
initial mem[412] = 16'he5c9;
initial mem[413] = 16'hec0a;
initial mem[414] = 16'hf28b;
initial mem[415] = 16'hf93a;
initial mem[416] = 16'h0;
initial mem[417] = 16'h641;
initial mem[418] = 16'hc70;
initial mem[419] = 16'h127b;
initial mem[420] = 16'h1852;
initial mem[421] = 16'h1deb;
initial mem[422] = 16'h233c;
initial mem[423] = 16'h283f;
initial mem[424] = 16'h2cf3;
initial mem[425] = 16'h3157;
initial mem[426] = 16'h356d;
initial mem[427] = 16'h3939;
initial mem[428] = 16'h3cbd;
initial mem[429] = 16'h3fff;
initial mem[430] = 16'h4303;
initial mem[431] = 16'h45ce;
initial mem[432] = 16'hb79b;
initial mem[433] = 16'hba32;
initial mem[434] = 16'hbcfd;
initial mem[435] = 16'hc001;
initial mem[436] = 16'hc343;
initial mem[437] = 16'hc6c7;
initial mem[438] = 16'hca93;
initial mem[439] = 16'hcea9;
initial mem[440] = 16'hd30d;
initial mem[441] = 16'hd7c1;
initial mem[442] = 16'hdcc4;
initial mem[443] = 16'he215;
initial mem[444] = 16'he7ae;
initial mem[445] = 16'hed85;
initial mem[446] = 16'hf390;
initial mem[447] = 16'hf9bf;
initial mem[448] = 16'h0;
initial mem[449] = 16'h5cf;
initial mem[450] = 16'hb8f;
initial mem[451] = 16'h1133;
initial mem[452] = 16'h16ad;
initial mem[453] = 16'h1bf3;
initial mem[454] = 16'h20fe;
initial mem[455] = 16'h25c7;
initial mem[456] = 16'h2a4d;
initial mem[457] = 16'h2e8e;
initial mem[458] = 16'h328a;
initial mem[459] = 16'h3644;
initial mem[460] = 16'h39be;
initial mem[461] = 16'h3cfb;
initial mem[462] = 16'h3fff;
initial mem[463] = 16'h42ce;
initial mem[464] = 16'hba94;
initial mem[465] = 16'hbd32;
initial mem[466] = 16'hc001;
initial mem[467] = 16'hc305;
initial mem[468] = 16'hc642;
initial mem[469] = 16'hc9bc;
initial mem[470] = 16'hcd76;
initial mem[471] = 16'hd172;
initial mem[472] = 16'hd5b3;
initial mem[473] = 16'hda39;
initial mem[474] = 16'hdf02;
initial mem[475] = 16'he40d;
initial mem[476] = 16'he953;
initial mem[477] = 16'heecd;
initial mem[478] = 16'hf471;
initial mem[479] = 16'hfa31;
initial mem[480] = 16'h0;
initial mem[481] = 16'h56c;
initial mem[482] = 16'hacd;
initial mem[483] = 16'h1015;
initial mem[484] = 16'h153c;
initial mem[485] = 16'h1a37;
initial mem[486] = 16'h1f01;
initial mem[487] = 16'h2394;
initial mem[488] = 16'h27ec;
initial mem[489] = 16'h2c09;
initial mem[490] = 16'h2fe9;
initial mem[491] = 16'h338f;
initial mem[492] = 16'h36fb;
initial mem[493] = 16'h3a30;
initial mem[494] = 16'h3d30;
initial mem[495] = 16'h3fff;
initial mem[496] = 16'hbd60;
initial mem[497] = 16'hc001;
initial mem[498] = 16'hc2d0;
initial mem[499] = 16'hc5d0;
initial mem[500] = 16'hc905;
initial mem[501] = 16'hcc71;
initial mem[502] = 16'hd017;
initial mem[503] = 16'hd3f7;
initial mem[504] = 16'hd814;
initial mem[505] = 16'hdc6c;
initial mem[506] = 16'he0ff;
initial mem[507] = 16'he5c9;
initial mem[508] = 16'heac4;
initial mem[509] = 16'hefeb;
initial mem[510] = 16'hf533;
initial mem[511] = 16'hfa94;
initial mem[512] = 16'hfffe;
initial mem[513] = 16'hfae7;
initial mem[514] = 16'hf5db;
initial mem[515] = 16'hf0e3;
initial mem[516] = 16'hec07;
initial mem[517] = 16'he74f;
initial mem[518] = 16'he2c2;
initial mem[519] = 16'hde63;
initial mem[520] = 16'hda36;
initial mem[521] = 16'hd63d;
initial mem[522] = 16'hd279;
initial mem[523] = 16'hceea;
initial mem[524] = 16'hcb8e;
initial mem[525] = 16'hc864;
initial mem[526] = 16'hc56b;
initial mem[527] = 16'hc29f;
initial mem[528] = 16'h4002;
initial mem[529] = 16'h3d61;
initial mem[530] = 16'h3a95;
initial mem[531] = 16'h379c;
initial mem[532] = 16'h3472;
initial mem[533] = 16'h3116;
initial mem[534] = 16'h2d87;
initial mem[535] = 16'h29c3;
initial mem[536] = 16'h25ca;
initial mem[537] = 16'h219d;
initial mem[538] = 16'h1d3e;
initial mem[539] = 16'h18b1;
initial mem[540] = 16'h13f9;
initial mem[541] = 16'hf1d;
initial mem[542] = 16'ha25;
initial mem[543] = 16'h519;
initial mem[544] = 16'hfffe;
initial mem[545] = 16'hfa91;
initial mem[546] = 16'hf530;
initial mem[547] = 16'hefe8;
initial mem[548] = 16'heac1;
initial mem[549] = 16'he5c6;
initial mem[550] = 16'he0fc;
initial mem[551] = 16'hdc69;
initial mem[552] = 16'hd811;
initial mem[553] = 16'hd3f4;
initial mem[554] = 16'hd014;
initial mem[555] = 16'hcc6e;
initial mem[556] = 16'hc902;
initial mem[557] = 16'hc5cd;
initial mem[558] = 16'hc2cd;
initial mem[559] = 16'hbffe;
initial mem[560] = 16'h42a3;
initial mem[561] = 16'h4002;
initial mem[562] = 16'h3d33;
initial mem[563] = 16'h3a33;
initial mem[564] = 16'h36fe;
initial mem[565] = 16'h3392;
initial mem[566] = 16'h2fec;
initial mem[567] = 16'h2c0c;
initial mem[568] = 16'h27ef;
initial mem[569] = 16'h2397;
initial mem[570] = 16'h1f04;
initial mem[571] = 16'h1a3a;
initial mem[572] = 16'h153f;
initial mem[573] = 16'h1018;
initial mem[574] = 16'had0;
initial mem[575] = 16'h56f;
initial mem[576] = 16'hfffe;
initial mem[577] = 16'hfa2e;
initial mem[578] = 16'hf46e;
initial mem[579] = 16'heeca;
initial mem[580] = 16'he950;
initial mem[581] = 16'he40a;
initial mem[582] = 16'hdeff;
initial mem[583] = 16'hda36;
initial mem[584] = 16'hd5b0;
initial mem[585] = 16'hd16f;
initial mem[586] = 16'hcd73;
initial mem[587] = 16'hc9b9;
initial mem[588] = 16'hc63f;
initial mem[589] = 16'hc302;
initial mem[590] = 16'hbffe;
initial mem[591] = 16'hbd2f;
initial mem[592] = 16'h456f;
initial mem[593] = 16'h42d1;
initial mem[594] = 16'h4002;
initial mem[595] = 16'h3cfe;
initial mem[596] = 16'h39c1;
initial mem[597] = 16'h3647;
initial mem[598] = 16'h328d;
initial mem[599] = 16'h2e91;
initial mem[600] = 16'h2a50;
initial mem[601] = 16'h25ca;
initial mem[602] = 16'h2101;
initial mem[603] = 16'h1bf6;
initial mem[604] = 16'h16b0;
initial mem[605] = 16'h1136;
initial mem[606] = 16'hb92;
initial mem[607] = 16'h5d2;
initial mem[608] = 16'hfffe;
initial mem[609] = 16'hf9bc;
initial mem[610] = 16'hf38d;
initial mem[611] = 16'hed82;
initial mem[612] = 16'he7ab;
initial mem[613] = 16'he212;
initial mem[614] = 16'hdcc1;
initial mem[615] = 16'hd7be;
initial mem[616] = 16'hd30a;
initial mem[617] = 16'hcea6;
initial mem[618] = 16'hca90;
initial mem[619] = 16'hc6c4;
initial mem[620] = 16'hc340;
initial mem[621] = 16'hbffe;
initial mem[622] = 16'hbcfa;
initial mem[623] = 16'hba2f;
initial mem[624] = 16'h4868;
initial mem[625] = 16'h45d1;
initial mem[626] = 16'h4306;
initial mem[627] = 16'h4002;
initial mem[628] = 16'h3cc0;
initial mem[629] = 16'h393c;
initial mem[630] = 16'h3570;
initial mem[631] = 16'h315a;
initial mem[632] = 16'h2cf6;
initial mem[633] = 16'h2842;
initial mem[634] = 16'h233f;
initial mem[635] = 16'h1dee;
initial mem[636] = 16'h1855;
initial mem[637] = 16'h127e;
initial mem[638] = 16'hc73;
initial mem[639] = 16'h644;
initial mem[640] = 16'hfffe;
initial mem[641] = 16'hf937;
initial mem[642] = 16'hf288;
initial mem[643] = 16'hec07;
initial mem[644] = 16'he5c6;
initial mem[645] = 16'hdfd2;
initial mem[646] = 16'hda36;
initial mem[647] = 16'hd4f6;
initial mem[648] = 16'hd014;
initial mem[649] = 16'hcb8e;
initial mem[650] = 16'hc761;
initial mem[651] = 16'hc388;
initial mem[652] = 16'hbffe;
initial mem[653] = 16'hbcbc;
initial mem[654] = 16'hb9bd;
initial mem[655] = 16'hb6fa;
initial mem[656] = 16'h4b92;
initial mem[657] = 16'h4906;
initial mem[658] = 16'h4643;
initial mem[659] = 16'h4344;
initial mem[660] = 16'h4002;
initial mem[661] = 16'h3c78;
initial mem[662] = 16'h389f;
initial mem[663] = 16'h3472;
initial mem[664] = 16'h2fec;
initial mem[665] = 16'h2b0a;
initial mem[666] = 16'h25ca;
initial mem[667] = 16'h202e;
initial mem[668] = 16'h1a3a;
initial mem[669] = 16'h13f9;
initial mem[670] = 16'hd78;
initial mem[671] = 16'h6c9;
initial mem[672] = 16'hfffe;
initial mem[673] = 16'hf89a;
initial mem[674] = 16'hf156;
initial mem[675] = 16'hea4b;
initial mem[676] = 16'he392;
initial mem[677] = 16'hdd3a;
initial mem[678] = 16'hd74d;
initial mem[679] = 16'hd1cf;
initial mem[680] = 16'hccc1;
initial mem[681] = 16'hc81d;
initial mem[682] = 16'hc3df;
initial mem[683] = 16'hbffe;
initial mem[684] = 16'hbc74;
initial mem[685] = 16'hb938;
initial mem[686] = 16'hb643;
initial mem[687] = 16'hb38e;
initial mem[688] = 16'h4eee;
initial mem[689] = 16'h4c72;
initial mem[690] = 16'h49bd;
initial mem[691] = 16'h46c8;
initial mem[692] = 16'h438c;
initial mem[693] = 16'h4002;
initial mem[694] = 16'h3c21;
initial mem[695] = 16'h37e3;
initial mem[696] = 16'h333f;
initial mem[697] = 16'h2e31;
initial mem[698] = 16'h28b3;
initial mem[699] = 16'h22c6;
initial mem[700] = 16'h1c6e;
initial mem[701] = 16'h15b5;
initial mem[702] = 16'heaa;
initial mem[703] = 16'h766;
initial mem[704] = 16'hfffe;
initial mem[705] = 16'hf7de;
initial mem[706] = 16'hefe8;
initial mem[707] = 16'he83e;
initial mem[708] = 16'he0fc;
initial mem[709] = 16'hda36;
initial mem[710] = 16'hd3f4;
initial mem[711] = 16'hce3a;
initial mem[712] = 16'hc902;
initial mem[713] = 16'hc447;
initial mem[714] = 16'hbffe;
initial mem[715] = 16'hbc1d;
initial mem[716] = 16'hb89b;
initial mem[717] = 16'hb56c;
initial mem[718] = 16'hb289;
initial mem[719] = 16'hafe8;
initial mem[720] = 16'h527d;
initial mem[721] = 16'h5018;
initial mem[722] = 16'h4d77;
initial mem[723] = 16'h4a94;
initial mem[724] = 16'h4765;
initial mem[725] = 16'h43e3;
initial mem[726] = 16'h4002;
initial mem[727] = 16'h3bb9;
initial mem[728] = 16'h36fe;
initial mem[729] = 16'h31c6;
initial mem[730] = 16'h2c0c;
initial mem[731] = 16'h25ca;
initial mem[732] = 16'h1f04;
initial mem[733] = 16'h17c2;
initial mem[734] = 16'h1018;
initial mem[735] = 16'h822;
initial mem[736] = 16'hfffe;
initial mem[737] = 16'hf6f9;
initial mem[738] = 16'hee2c;
initial mem[739] = 16'he5c6;
initial mem[740] = 16'hdde9;
initial mem[741] = 16'hd6ab;
initial mem[742] = 16'hd014;
initial mem[743] = 16'hca20;
initial mem[744] = 16'hc4c8;
initial mem[745] = 16'hbffe;
initial mem[746] = 16'hbbb5;
initial mem[747] = 16'hb7df;
initial mem[748] = 16'hb46e;
initial mem[749] = 16'hb156;
initial mem[750] = 16'hae8d;
initial mem[751] = 16'hac08;
initial mem[752] = 16'h5641;
initial mem[753] = 16'h53f8;
initial mem[754] = 16'h5173;
initial mem[755] = 16'h4eaa;
initial mem[756] = 16'h4b92;
initial mem[757] = 16'h4821;
initial mem[758] = 16'h444b;
initial mem[759] = 16'h4002;
initial mem[760] = 16'h3b38;
initial mem[761] = 16'h35e0;
initial mem[762] = 16'h2fec;
initial mem[763] = 16'h2955;
initial mem[764] = 16'h2217;
initial mem[765] = 16'h1a3a;
initial mem[766] = 16'h11d4;
initial mem[767] = 16'h907;
initial mem[768] = 16'hfffe;
initial mem[769] = 16'hf5db;
initial mem[770] = 16'hec07;
initial mem[771] = 16'he2c2;
initial mem[772] = 16'hda36;
initial mem[773] = 16'hd279;
initial mem[774] = 16'hcb8e;
initial mem[775] = 16'hc56b;
initial mem[776] = 16'hbffe;
initial mem[777] = 16'hbb34;
initial mem[778] = 16'hb6fa;
initial mem[779] = 16'hb33b;
initial mem[780] = 16'hafe8;
initial mem[781] = 16'hacf2;
initial mem[782] = 16'haa4c;
initial mem[783] = 16'ha7eb;
initial mem[784] = 16'h5a3a;
initial mem[785] = 16'h5815;
initial mem[786] = 16'h55b4;
initial mem[787] = 16'h530e;
initial mem[788] = 16'h5018;
initial mem[789] = 16'h4cc5;
initial mem[790] = 16'h4906;
initial mem[791] = 16'h44cc;
initial mem[792] = 16'h4002;
initial mem[793] = 16'h3a95;
initial mem[794] = 16'h3472;
initial mem[795] = 16'h2d87;
initial mem[796] = 16'h25ca;
initial mem[797] = 16'h1d3e;
initial mem[798] = 16'h13f9;
initial mem[799] = 16'ha25;
initial mem[800] = 16'hfffe;
initial mem[801] = 16'hf46e;
initial mem[802] = 16'he950;
initial mem[803] = 16'hdeff;
initial mem[804] = 16'hd5b0;
initial mem[805] = 16'hcd73;
initial mem[806] = 16'hc63f;
initial mem[807] = 16'hbffe;
initial mem[808] = 16'hba91;
initial mem[809] = 16'hb5dc;
initial mem[810] = 16'hb1c2;
initial mem[811] = 16'hae2d;
initial mem[812] = 16'hab06;
initial mem[813] = 16'ha83e;
initial mem[814] = 16'ha5c6;
initial mem[815] = 16'ha393;
initial mem[816] = 16'h5e67;
initial mem[817] = 16'h5c6d;
initial mem[818] = 16'h5a3a;
initial mem[819] = 16'h57c2;
initial mem[820] = 16'h54fa;
initial mem[821] = 16'h51d3;
initial mem[822] = 16'h4e3e;
initial mem[823] = 16'h4a24;
initial mem[824] = 16'h456f;
initial mem[825] = 16'h4002;
initial mem[826] = 16'h39c1;
initial mem[827] = 16'h328d;
initial mem[828] = 16'h2a50;
initial mem[829] = 16'h2101;
initial mem[830] = 16'h16b0;
initial mem[831] = 16'hb92;
initial mem[832] = 16'hfffe;
initial mem[833] = 16'hf288;
initial mem[834] = 16'he5c6;
initial mem[835] = 16'hda36;
initial mem[836] = 16'hd014;
initial mem[837] = 16'hc761;
initial mem[838] = 16'hbffe;
initial mem[839] = 16'hb9bd;
initial mem[840] = 16'hb46e;
initial mem[841] = 16'hafe8;
initial mem[842] = 16'hac08;
initial mem[843] = 16'ha8af;
initial mem[844] = 16'ha5c6;
initial mem[845] = 16'ha33b;
initial mem[846] = 16'ha0fd;
initial mem[847] = 16'h9f00;
initial mem[848] = 16'h62c6;
initial mem[849] = 16'h6100;
initial mem[850] = 16'h5f03;
initial mem[851] = 16'h5cc5;
initial mem[852] = 16'h5a3a;
initial mem[853] = 16'h5751;
initial mem[854] = 16'h53f8;
initial mem[855] = 16'h5018;
initial mem[856] = 16'h4b92;
initial mem[857] = 16'h4643;
initial mem[858] = 16'h4002;
initial mem[859] = 16'h389f;
initial mem[860] = 16'h2fec;
initial mem[861] = 16'h25ca;
initial mem[862] = 16'h1a3a;
initial mem[863] = 16'hd78;
initial mem[864] = 16'hfffe;
initial mem[865] = 16'hefe8;
initial mem[866] = 16'he0fc;
initial mem[867] = 16'hd3f4;
initial mem[868] = 16'hc902;
initial mem[869] = 16'hbffe;
initial mem[870] = 16'hb89b;
initial mem[871] = 16'hb289;
initial mem[872] = 16'had83;
initial mem[873] = 16'ha951;
initial mem[874] = 16'ha5c6;
initial mem[875] = 16'ha2c2;
initial mem[876] = 16'ha02a;
initial mem[877] = 16'h9dea;
initial mem[878] = 16'h9bf2;
initial mem[879] = 16'h9a36;
initial mem[880] = 16'h6753;
initial mem[881] = 16'h65ca;
initial mem[882] = 16'h640e;
initial mem[883] = 16'h6216;
initial mem[884] = 16'h5fd6;
initial mem[885] = 16'h5d3e;
initial mem[886] = 16'h5a3a;
initial mem[887] = 16'h56af;
initial mem[888] = 16'h527d;
initial mem[889] = 16'h4d77;
initial mem[890] = 16'h4765;
initial mem[891] = 16'h4002;
initial mem[892] = 16'h36fe;
initial mem[893] = 16'h2c0c;
initial mem[894] = 16'h1f04;
initial mem[895] = 16'h1018;
initial mem[896] = 16'hfffe;
initial mem[897] = 16'hec07;
initial mem[898] = 16'hda36;
initial mem[899] = 16'hcb8e;
initial mem[900] = 16'hbffe;
initial mem[901] = 16'hb6fa;
initial mem[902] = 16'hafe8;
initial mem[903] = 16'haa4c;
initial mem[904] = 16'ha5c6;
initial mem[905] = 16'ha213;
initial mem[906] = 16'h9f00;
initial mem[907] = 16'h9c6a;
initial mem[908] = 16'h9a36;
initial mem[909] = 16'h9851;
initial mem[910] = 16'h96ac;
initial mem[911] = 16'h953b;
initial mem[912] = 16'h6c0b;
initial mem[913] = 16'h6ac5;
initial mem[914] = 16'h6954;
initial mem[915] = 16'h67af;
initial mem[916] = 16'h65ca;
initial mem[917] = 16'h6396;
initial mem[918] = 16'h6100;
initial mem[919] = 16'h5ded;
initial mem[920] = 16'h5a3a;
initial mem[921] = 16'h55b4;
initial mem[922] = 16'h5018;
initial mem[923] = 16'h4906;
initial mem[924] = 16'h4002;
initial mem[925] = 16'h3472;
initial mem[926] = 16'h25ca;
initial mem[927] = 16'h13f9;
initial mem[928] = 16'hfffe;
initial mem[929] = 16'he5c6;
initial mem[930] = 16'hd014;
initial mem[931] = 16'hbffe;
initial mem[932] = 16'hb46e;
initial mem[933] = 16'hac08;
initial mem[934] = 16'ha5c6;
initial mem[935] = 16'ha0fd;
initial mem[936] = 16'h9d3a;
initial mem[937] = 16'h9a36;
initial mem[938] = 16'h97be;
initial mem[939] = 16'h95b1;
initial mem[940] = 16'h93f5;
initial mem[941] = 16'h927a;
initial mem[942] = 16'h9132;
initial mem[943] = 16'h9014;
initial mem[944] = 16'h70e7;
initial mem[945] = 16'h6fec;
initial mem[946] = 16'h6ece;
initial mem[947] = 16'h6d86;
initial mem[948] = 16'h6c0b;
initial mem[949] = 16'h6a4f;
initial mem[950] = 16'h6842;
initial mem[951] = 16'h65ca;
initial mem[952] = 16'h62c6;
initial mem[953] = 16'h5f03;
initial mem[954] = 16'h5a3a;
initial mem[955] = 16'h53f8;
initial mem[956] = 16'h4b92;
initial mem[957] = 16'h4002;
initial mem[958] = 16'h2fec;
initial mem[959] = 16'h1a3a;
initial mem[960] = 16'hfffe;
initial mem[961] = 16'hda36;
initial mem[962] = 16'hbffe;
initial mem[963] = 16'hafe8;
initial mem[964] = 16'ha5c6;
initial mem[965] = 16'h9f00;
initial mem[966] = 16'h9a36;
initial mem[967] = 16'h96ac;
initial mem[968] = 16'h93f5;
initial mem[969] = 16'h91d0;
initial mem[970] = 16'h9014;
initial mem[971] = 16'h8ea6;
initial mem[972] = 16'h8d74;
initial mem[973] = 16'h8c6f;
initial mem[974] = 16'h8b8e;
initial mem[975] = 16'h8acc;
initial mem[976] = 16'h75df;
initial mem[977] = 16'h7534;
initial mem[978] = 16'h7472;
initial mem[979] = 16'h7391;
initial mem[980] = 16'h728c;
initial mem[981] = 16'h715a;
initial mem[982] = 16'h6fec;
initial mem[983] = 16'h6e30;
initial mem[984] = 16'h6c0b;
initial mem[985] = 16'h6954;
initial mem[986] = 16'h65ca;
initial mem[987] = 16'h6100;
initial mem[988] = 16'h5a3a;
initial mem[989] = 16'h5018;
initial mem[990] = 16'h4002;
initial mem[991] = 16'h25ca;
initial mem[992] = 16'hfffe;
initial mem[993] = 16'hbffe;
initial mem[994] = 16'ha5c6;
initial mem[995] = 16'h9a36;
initial mem[996] = 16'h93f5;
initial mem[997] = 16'h9014;
initial mem[998] = 16'h8d74;
initial mem[999] = 16'h8b8e;
initial mem[1000] = 16'h8a21;
initial mem[1001] = 16'h8903;
initial mem[1002] = 16'h881e;
initial mem[1003] = 16'h8762;
initial mem[1004] = 16'h86c5;
initial mem[1005] = 16'h8640;
initial mem[1006] = 16'h85ce;
initial mem[1007] = 16'h856b;
initial mem[1008] = 16'h7aeb;
initial mem[1009] = 16'h7a95;
initial mem[1010] = 16'h7a32;
initial mem[1011] = 16'h79c0;
initial mem[1012] = 16'h793b;
initial mem[1013] = 16'h789e;
initial mem[1014] = 16'h77e2;
initial mem[1015] = 16'h76fd;
initial mem[1016] = 16'h75df;
initial mem[1017] = 16'h7472;
initial mem[1018] = 16'h728c;
initial mem[1019] = 16'h6fec;
initial mem[1020] = 16'h6c0b;
initial mem[1021] = 16'h65ca;
initial mem[1022] = 16'h5a3a;
initial mem[1023] = 16'h4002;
always @(posedge clk) begin
	data <= mem[addr];
end
endmodule
