module argTable(input clk, input [9:0] addr, output reg [15:0] data);
reg [15:0] mem [0:1023];
initial mem[0] = 16'h0;
initial mem[1] = 16'h7fff;
initial mem[2] = 16'h7fff;
initial mem[3] = 16'h7fff;
initial mem[4] = 16'h7fff;
initial mem[5] = 16'h7fff;
initial mem[6] = 16'h7fff;
initial mem[7] = 16'h7fff;
initial mem[8] = 16'h7fff;
initial mem[9] = 16'h7fff;
initial mem[10] = 16'h7fff;
initial mem[11] = 16'h7fff;
initial mem[12] = 16'h7fff;
initial mem[13] = 16'h7fff;
initial mem[14] = 16'h7fff;
initial mem[15] = 16'h7fff;
initial mem[16] = 16'h8001;
initial mem[17] = 16'h8001;
initial mem[18] = 16'h8001;
initial mem[19] = 16'h8001;
initial mem[20] = 16'h8001;
initial mem[21] = 16'h8001;
initial mem[22] = 16'h8001;
initial mem[23] = 16'h8001;
initial mem[24] = 16'h8001;
initial mem[25] = 16'h8001;
initial mem[26] = 16'h8001;
initial mem[27] = 16'h8001;
initial mem[28] = 16'h8001;
initial mem[29] = 16'h8001;
initial mem[30] = 16'h8001;
initial mem[31] = 16'h8001;
initial mem[32] = 16'h0;
initial mem[33] = 16'h3fff;
initial mem[34] = 16'h5a37;
initial mem[35] = 16'h65c7;
initial mem[36] = 16'h6c08;
initial mem[37] = 16'h6fe9;
initial mem[38] = 16'h7289;
initial mem[39] = 16'h746f;
initial mem[40] = 16'h75dc;
initial mem[41] = 16'h76fa;
initial mem[42] = 16'h77df;
initial mem[43] = 16'h789b;
initial mem[44] = 16'h7938;
initial mem[45] = 16'h79bd;
initial mem[46] = 16'h7a2f;
initial mem[47] = 16'h7a92;
initial mem[48] = 16'h8518;
initial mem[49] = 16'h856e;
initial mem[50] = 16'h85d1;
initial mem[51] = 16'h8643;
initial mem[52] = 16'h86c8;
initial mem[53] = 16'h8765;
initial mem[54] = 16'h8821;
initial mem[55] = 16'h8906;
initial mem[56] = 16'h8a24;
initial mem[57] = 16'h8b91;
initial mem[58] = 16'h8d77;
initial mem[59] = 16'h9017;
initial mem[60] = 16'h93f8;
initial mem[61] = 16'h9a39;
initial mem[62] = 16'ha5c9;
initial mem[63] = 16'hc001;
initial mem[64] = 16'h0;
initial mem[65] = 16'h7fff;
initial mem[66] = 16'h7fff;
initial mem[67] = 16'h7fff;
initial mem[68] = 16'h7fff;
initial mem[69] = 16'h7fff;
initial mem[70] = 16'h7fff;
initial mem[71] = 16'h7fff;
initial mem[72] = 16'h7fff;
initial mem[73] = 16'h7fff;
initial mem[74] = 16'h7fff;
initial mem[75] = 16'h7fff;
initial mem[76] = 16'h7fff;
initial mem[77] = 16'h7fff;
initial mem[78] = 16'h7fff;
initial mem[79] = 16'h7fff;
initial mem[80] = 16'h8001;
initial mem[81] = 16'h8001;
initial mem[82] = 16'h8001;
initial mem[83] = 16'h8001;
initial mem[84] = 16'h8001;
initial mem[85] = 16'h8001;
initial mem[86] = 16'h8001;
initial mem[87] = 16'h8001;
initial mem[88] = 16'h8001;
initial mem[89] = 16'h8001;
initial mem[90] = 16'h8001;
initial mem[91] = 16'h8001;
initial mem[92] = 16'h8001;
initial mem[93] = 16'h8001;
initial mem[94] = 16'h8001;
initial mem[95] = 16'h8001;
initial mem[96] = 16'h0;
initial mem[97] = 16'h3fff;
initial mem[98] = 16'h5a37;
initial mem[99] = 16'h65c7;
initial mem[100] = 16'h6c08;
initial mem[101] = 16'h6fe9;
initial mem[102] = 16'h7289;
initial mem[103] = 16'h746f;
initial mem[104] = 16'h75dc;
initial mem[105] = 16'h76fa;
initial mem[106] = 16'h77df;
initial mem[107] = 16'h789b;
initial mem[108] = 16'h7938;
initial mem[109] = 16'h79bd;
initial mem[110] = 16'h7a2f;
initial mem[111] = 16'h7a92;
initial mem[112] = 16'h8518;
initial mem[113] = 16'h856e;
initial mem[114] = 16'h85d1;
initial mem[115] = 16'h8643;
initial mem[116] = 16'h86c8;
initial mem[117] = 16'h8765;
initial mem[118] = 16'h8821;
initial mem[119] = 16'h8906;
initial mem[120] = 16'h8a24;
initial mem[121] = 16'h8b91;
initial mem[122] = 16'h8d77;
initial mem[123] = 16'h9017;
initial mem[124] = 16'h93f8;
initial mem[125] = 16'h9a39;
initial mem[126] = 16'ha5c9;
initial mem[127] = 16'hc001;
initial mem[128] = 16'h0;
initial mem[129] = 16'h7fff;
initial mem[130] = 16'h7fff;
initial mem[131] = 16'h7fff;
initial mem[132] = 16'h7fff;
initial mem[133] = 16'h7fff;
initial mem[134] = 16'h7fff;
initial mem[135] = 16'h7fff;
initial mem[136] = 16'h7fff;
initial mem[137] = 16'h7fff;
initial mem[138] = 16'h7fff;
initial mem[139] = 16'h7fff;
initial mem[140] = 16'h7fff;
initial mem[141] = 16'h7fff;
initial mem[142] = 16'h7fff;
initial mem[143] = 16'h7fff;
initial mem[144] = 16'h8001;
initial mem[145] = 16'h8001;
initial mem[146] = 16'h8001;
initial mem[147] = 16'h8001;
initial mem[148] = 16'h8001;
initial mem[149] = 16'h8001;
initial mem[150] = 16'h8001;
initial mem[151] = 16'h8001;
initial mem[152] = 16'h8001;
initial mem[153] = 16'h8001;
initial mem[154] = 16'h8001;
initial mem[155] = 16'h8001;
initial mem[156] = 16'h8001;
initial mem[157] = 16'h8001;
initial mem[158] = 16'h8001;
initial mem[159] = 16'h8001;
initial mem[160] = 16'h0;
initial mem[161] = 16'h3fff;
initial mem[162] = 16'h5a37;
initial mem[163] = 16'h65c7;
initial mem[164] = 16'h6c08;
initial mem[165] = 16'h6fe9;
initial mem[166] = 16'h7289;
initial mem[167] = 16'h746f;
initial mem[168] = 16'h75dc;
initial mem[169] = 16'h76fa;
initial mem[170] = 16'h77df;
initial mem[171] = 16'h789b;
initial mem[172] = 16'h7938;
initial mem[173] = 16'h79bd;
initial mem[174] = 16'h7a2f;
initial mem[175] = 16'h7a92;
initial mem[176] = 16'h8518;
initial mem[177] = 16'h856e;
initial mem[178] = 16'h85d1;
initial mem[179] = 16'h8643;
initial mem[180] = 16'h86c8;
initial mem[181] = 16'h8765;
initial mem[182] = 16'h8821;
initial mem[183] = 16'h8906;
initial mem[184] = 16'h8a24;
initial mem[185] = 16'h8b91;
initial mem[186] = 16'h8d77;
initial mem[187] = 16'h9017;
initial mem[188] = 16'h93f8;
initial mem[189] = 16'h9a39;
initial mem[190] = 16'ha5c9;
initial mem[191] = 16'hc001;
initial mem[192] = 16'h0;
initial mem[193] = 16'h7fff;
initial mem[194] = 16'h7fff;
initial mem[195] = 16'h7fff;
initial mem[196] = 16'h7fff;
initial mem[197] = 16'h7fff;
initial mem[198] = 16'h7fff;
initial mem[199] = 16'h7fff;
initial mem[200] = 16'h7fff;
initial mem[201] = 16'h7fff;
initial mem[202] = 16'h7fff;
initial mem[203] = 16'h7fff;
initial mem[204] = 16'h7fff;
initial mem[205] = 16'h7fff;
initial mem[206] = 16'h7fff;
initial mem[207] = 16'h7fff;
initial mem[208] = 16'h8001;
initial mem[209] = 16'h8001;
initial mem[210] = 16'h8001;
initial mem[211] = 16'h8001;
initial mem[212] = 16'h8001;
initial mem[213] = 16'h8001;
initial mem[214] = 16'h8001;
initial mem[215] = 16'h8001;
initial mem[216] = 16'h8001;
initial mem[217] = 16'h8001;
initial mem[218] = 16'h8001;
initial mem[219] = 16'h8001;
initial mem[220] = 16'h8001;
initial mem[221] = 16'h8001;
initial mem[222] = 16'h8001;
initial mem[223] = 16'h8001;
initial mem[224] = 16'h0;
initial mem[225] = 16'h3fff;
initial mem[226] = 16'h5a37;
initial mem[227] = 16'h65c7;
initial mem[228] = 16'h6c08;
initial mem[229] = 16'h6fe9;
initial mem[230] = 16'h7289;
initial mem[231] = 16'h746f;
initial mem[232] = 16'h75dc;
initial mem[233] = 16'h76fa;
initial mem[234] = 16'h77df;
initial mem[235] = 16'h789b;
initial mem[236] = 16'h7938;
initial mem[237] = 16'h79bd;
initial mem[238] = 16'h7a2f;
initial mem[239] = 16'h7a92;
initial mem[240] = 16'h8518;
initial mem[241] = 16'h856e;
initial mem[242] = 16'h85d1;
initial mem[243] = 16'h8643;
initial mem[244] = 16'h86c8;
initial mem[245] = 16'h8765;
initial mem[246] = 16'h8821;
initial mem[247] = 16'h8906;
initial mem[248] = 16'h8a24;
initial mem[249] = 16'h8b91;
initial mem[250] = 16'h8d77;
initial mem[251] = 16'h9017;
initial mem[252] = 16'h93f8;
initial mem[253] = 16'h9a39;
initial mem[254] = 16'ha5c9;
initial mem[255] = 16'hc001;
initial mem[256] = 16'h0;
initial mem[257] = 16'h7fff;
initial mem[258] = 16'h7fff;
initial mem[259] = 16'h7fff;
initial mem[260] = 16'h7fff;
initial mem[261] = 16'h7fff;
initial mem[262] = 16'h7fff;
initial mem[263] = 16'h7fff;
initial mem[264] = 16'h7fff;
initial mem[265] = 16'h7fff;
initial mem[266] = 16'h7fff;
initial mem[267] = 16'h7fff;
initial mem[268] = 16'h7fff;
initial mem[269] = 16'h7fff;
initial mem[270] = 16'h7fff;
initial mem[271] = 16'h7fff;
initial mem[272] = 16'h8001;
initial mem[273] = 16'h8001;
initial mem[274] = 16'h8001;
initial mem[275] = 16'h8001;
initial mem[276] = 16'h8001;
initial mem[277] = 16'h8001;
initial mem[278] = 16'h8001;
initial mem[279] = 16'h8001;
initial mem[280] = 16'h8001;
initial mem[281] = 16'h8001;
initial mem[282] = 16'h8001;
initial mem[283] = 16'h8001;
initial mem[284] = 16'h8001;
initial mem[285] = 16'h8001;
initial mem[286] = 16'h8001;
initial mem[287] = 16'h8001;
initial mem[288] = 16'h0;
initial mem[289] = 16'h3fff;
initial mem[290] = 16'h5a37;
initial mem[291] = 16'h65c7;
initial mem[292] = 16'h6c08;
initial mem[293] = 16'h6fe9;
initial mem[294] = 16'h7289;
initial mem[295] = 16'h746f;
initial mem[296] = 16'h75dc;
initial mem[297] = 16'h76fa;
initial mem[298] = 16'h77df;
initial mem[299] = 16'h789b;
initial mem[300] = 16'h7938;
initial mem[301] = 16'h79bd;
initial mem[302] = 16'h7a2f;
initial mem[303] = 16'h7a92;
initial mem[304] = 16'h8518;
initial mem[305] = 16'h856e;
initial mem[306] = 16'h85d1;
initial mem[307] = 16'h8643;
initial mem[308] = 16'h86c8;
initial mem[309] = 16'h8765;
initial mem[310] = 16'h8821;
initial mem[311] = 16'h8906;
initial mem[312] = 16'h8a24;
initial mem[313] = 16'h8b91;
initial mem[314] = 16'h8d77;
initial mem[315] = 16'h9017;
initial mem[316] = 16'h93f8;
initial mem[317] = 16'h9a39;
initial mem[318] = 16'ha5c9;
initial mem[319] = 16'hc001;
initial mem[320] = 16'h0;
initial mem[321] = 16'h7fff;
initial mem[322] = 16'h7fff;
initial mem[323] = 16'h7fff;
initial mem[324] = 16'h7fff;
initial mem[325] = 16'h7fff;
initial mem[326] = 16'h7fff;
initial mem[327] = 16'h7fff;
initial mem[328] = 16'h7fff;
initial mem[329] = 16'h7fff;
initial mem[330] = 16'h7fff;
initial mem[331] = 16'h7fff;
initial mem[332] = 16'h7fff;
initial mem[333] = 16'h7fff;
initial mem[334] = 16'h7fff;
initial mem[335] = 16'h7fff;
initial mem[336] = 16'h8001;
initial mem[337] = 16'h8001;
initial mem[338] = 16'h8001;
initial mem[339] = 16'h8001;
initial mem[340] = 16'h8001;
initial mem[341] = 16'h8001;
initial mem[342] = 16'h8001;
initial mem[343] = 16'h8001;
initial mem[344] = 16'h8001;
initial mem[345] = 16'h8001;
initial mem[346] = 16'h8001;
initial mem[347] = 16'h8001;
initial mem[348] = 16'h8001;
initial mem[349] = 16'h8001;
initial mem[350] = 16'h8001;
initial mem[351] = 16'h8001;
initial mem[352] = 16'h0;
initial mem[353] = 16'h3fff;
initial mem[354] = 16'h5a37;
initial mem[355] = 16'h65c7;
initial mem[356] = 16'h6c08;
initial mem[357] = 16'h6fe9;
initial mem[358] = 16'h7289;
initial mem[359] = 16'h746f;
initial mem[360] = 16'h75dc;
initial mem[361] = 16'h76fa;
initial mem[362] = 16'h77df;
initial mem[363] = 16'h789b;
initial mem[364] = 16'h7938;
initial mem[365] = 16'h79bd;
initial mem[366] = 16'h7a2f;
initial mem[367] = 16'h7a92;
initial mem[368] = 16'h8518;
initial mem[369] = 16'h856e;
initial mem[370] = 16'h85d1;
initial mem[371] = 16'h8643;
initial mem[372] = 16'h86c8;
initial mem[373] = 16'h8765;
initial mem[374] = 16'h8821;
initial mem[375] = 16'h8906;
initial mem[376] = 16'h8a24;
initial mem[377] = 16'h8b91;
initial mem[378] = 16'h8d77;
initial mem[379] = 16'h9017;
initial mem[380] = 16'h93f8;
initial mem[381] = 16'h9a39;
initial mem[382] = 16'ha5c9;
initial mem[383] = 16'hc001;
initial mem[384] = 16'h0;
initial mem[385] = 16'h7fff;
initial mem[386] = 16'h7fff;
initial mem[387] = 16'h7fff;
initial mem[388] = 16'h7fff;
initial mem[389] = 16'h7fff;
initial mem[390] = 16'h7fff;
initial mem[391] = 16'h7fff;
initial mem[392] = 16'h7fff;
initial mem[393] = 16'h7fff;
initial mem[394] = 16'h7fff;
initial mem[395] = 16'h7fff;
initial mem[396] = 16'h7fff;
initial mem[397] = 16'h7fff;
initial mem[398] = 16'h7fff;
initial mem[399] = 16'h7fff;
initial mem[400] = 16'h8001;
initial mem[401] = 16'h8001;
initial mem[402] = 16'h8001;
initial mem[403] = 16'h8001;
initial mem[404] = 16'h8001;
initial mem[405] = 16'h8001;
initial mem[406] = 16'h8001;
initial mem[407] = 16'h8001;
initial mem[408] = 16'h8001;
initial mem[409] = 16'h8001;
initial mem[410] = 16'h8001;
initial mem[411] = 16'h8001;
initial mem[412] = 16'h8001;
initial mem[413] = 16'h8001;
initial mem[414] = 16'h8001;
initial mem[415] = 16'h8001;
initial mem[416] = 16'h0;
initial mem[417] = 16'h3fff;
initial mem[418] = 16'h5a37;
initial mem[419] = 16'h65c7;
initial mem[420] = 16'h6c08;
initial mem[421] = 16'h6fe9;
initial mem[422] = 16'h7289;
initial mem[423] = 16'h746f;
initial mem[424] = 16'h75dc;
initial mem[425] = 16'h76fa;
initial mem[426] = 16'h77df;
initial mem[427] = 16'h789b;
initial mem[428] = 16'h7938;
initial mem[429] = 16'h79bd;
initial mem[430] = 16'h7a2f;
initial mem[431] = 16'h7a92;
initial mem[432] = 16'h8518;
initial mem[433] = 16'h856e;
initial mem[434] = 16'h85d1;
initial mem[435] = 16'h8643;
initial mem[436] = 16'h86c8;
initial mem[437] = 16'h8765;
initial mem[438] = 16'h8821;
initial mem[439] = 16'h8906;
initial mem[440] = 16'h8a24;
initial mem[441] = 16'h8b91;
initial mem[442] = 16'h8d77;
initial mem[443] = 16'h9017;
initial mem[444] = 16'h93f8;
initial mem[445] = 16'h9a39;
initial mem[446] = 16'ha5c9;
initial mem[447] = 16'hc001;
initial mem[448] = 16'h0;
initial mem[449] = 16'h7fff;
initial mem[450] = 16'h7fff;
initial mem[451] = 16'h7fff;
initial mem[452] = 16'h7fff;
initial mem[453] = 16'h7fff;
initial mem[454] = 16'h7fff;
initial mem[455] = 16'h7fff;
initial mem[456] = 16'h7fff;
initial mem[457] = 16'h7fff;
initial mem[458] = 16'h7fff;
initial mem[459] = 16'h7fff;
initial mem[460] = 16'h7fff;
initial mem[461] = 16'h7fff;
initial mem[462] = 16'h7fff;
initial mem[463] = 16'h7fff;
initial mem[464] = 16'h8001;
initial mem[465] = 16'h8001;
initial mem[466] = 16'h8001;
initial mem[467] = 16'h8001;
initial mem[468] = 16'h8001;
initial mem[469] = 16'h8001;
initial mem[470] = 16'h8001;
initial mem[471] = 16'h8001;
initial mem[472] = 16'h8001;
initial mem[473] = 16'h8001;
initial mem[474] = 16'h8001;
initial mem[475] = 16'h8001;
initial mem[476] = 16'h8001;
initial mem[477] = 16'h8001;
initial mem[478] = 16'h8001;
initial mem[479] = 16'h8001;
initial mem[480] = 16'h0;
initial mem[481] = 16'h3fff;
initial mem[482] = 16'h5a37;
initial mem[483] = 16'h65c7;
initial mem[484] = 16'h6c08;
initial mem[485] = 16'h6fe9;
initial mem[486] = 16'h7289;
initial mem[487] = 16'h746f;
initial mem[488] = 16'h75dc;
initial mem[489] = 16'h76fa;
initial mem[490] = 16'h77df;
initial mem[491] = 16'h789b;
initial mem[492] = 16'h7938;
initial mem[493] = 16'h79bd;
initial mem[494] = 16'h7a2f;
initial mem[495] = 16'h7a92;
initial mem[496] = 16'h8518;
initial mem[497] = 16'h856e;
initial mem[498] = 16'h85d1;
initial mem[499] = 16'h8643;
initial mem[500] = 16'h86c8;
initial mem[501] = 16'h8765;
initial mem[502] = 16'h8821;
initial mem[503] = 16'h8906;
initial mem[504] = 16'h8a24;
initial mem[505] = 16'h8b91;
initial mem[506] = 16'h8d77;
initial mem[507] = 16'h9017;
initial mem[508] = 16'h93f8;
initial mem[509] = 16'h9a39;
initial mem[510] = 16'ha5c9;
initial mem[511] = 16'hc001;
initial mem[512] = 16'h0;
initial mem[513] = 16'h7fff;
initial mem[514] = 16'h7fff;
initial mem[515] = 16'h7fff;
initial mem[516] = 16'h7fff;
initial mem[517] = 16'h7fff;
initial mem[518] = 16'h7fff;
initial mem[519] = 16'h7fff;
initial mem[520] = 16'h7fff;
initial mem[521] = 16'h7fff;
initial mem[522] = 16'h7fff;
initial mem[523] = 16'h7fff;
initial mem[524] = 16'h7fff;
initial mem[525] = 16'h7fff;
initial mem[526] = 16'h7fff;
initial mem[527] = 16'h7fff;
initial mem[528] = 16'h8001;
initial mem[529] = 16'h8001;
initial mem[530] = 16'h8001;
initial mem[531] = 16'h8001;
initial mem[532] = 16'h8001;
initial mem[533] = 16'h8001;
initial mem[534] = 16'h8001;
initial mem[535] = 16'h8001;
initial mem[536] = 16'h8001;
initial mem[537] = 16'h8001;
initial mem[538] = 16'h8001;
initial mem[539] = 16'h8001;
initial mem[540] = 16'h8001;
initial mem[541] = 16'h8001;
initial mem[542] = 16'h8001;
initial mem[543] = 16'h8001;
initial mem[544] = 16'h0;
initial mem[545] = 16'h3fff;
initial mem[546] = 16'h5a37;
initial mem[547] = 16'h65c7;
initial mem[548] = 16'h6c08;
initial mem[549] = 16'h6fe9;
initial mem[550] = 16'h7289;
initial mem[551] = 16'h746f;
initial mem[552] = 16'h75dc;
initial mem[553] = 16'h76fa;
initial mem[554] = 16'h77df;
initial mem[555] = 16'h789b;
initial mem[556] = 16'h7938;
initial mem[557] = 16'h79bd;
initial mem[558] = 16'h7a2f;
initial mem[559] = 16'h7a92;
initial mem[560] = 16'h8518;
initial mem[561] = 16'h856e;
initial mem[562] = 16'h85d1;
initial mem[563] = 16'h8643;
initial mem[564] = 16'h86c8;
initial mem[565] = 16'h8765;
initial mem[566] = 16'h8821;
initial mem[567] = 16'h8906;
initial mem[568] = 16'h8a24;
initial mem[569] = 16'h8b91;
initial mem[570] = 16'h8d77;
initial mem[571] = 16'h9017;
initial mem[572] = 16'h93f8;
initial mem[573] = 16'h9a39;
initial mem[574] = 16'ha5c9;
initial mem[575] = 16'hc001;
initial mem[576] = 16'h0;
initial mem[577] = 16'h7fff;
initial mem[578] = 16'h7fff;
initial mem[579] = 16'h7fff;
initial mem[580] = 16'h7fff;
initial mem[581] = 16'h7fff;
initial mem[582] = 16'h7fff;
initial mem[583] = 16'h7fff;
initial mem[584] = 16'h7fff;
initial mem[585] = 16'h7fff;
initial mem[586] = 16'h7fff;
initial mem[587] = 16'h7fff;
initial mem[588] = 16'h7fff;
initial mem[589] = 16'h7fff;
initial mem[590] = 16'h7fff;
initial mem[591] = 16'h7fff;
initial mem[592] = 16'h8001;
initial mem[593] = 16'h8001;
initial mem[594] = 16'h8001;
initial mem[595] = 16'h8001;
initial mem[596] = 16'h8001;
initial mem[597] = 16'h8001;
initial mem[598] = 16'h8001;
initial mem[599] = 16'h8001;
initial mem[600] = 16'h8001;
initial mem[601] = 16'h8001;
initial mem[602] = 16'h8001;
initial mem[603] = 16'h8001;
initial mem[604] = 16'h8001;
initial mem[605] = 16'h8001;
initial mem[606] = 16'h8001;
initial mem[607] = 16'h8001;
initial mem[608] = 16'h0;
initial mem[609] = 16'h3fff;
initial mem[610] = 16'h5a37;
initial mem[611] = 16'h65c7;
initial mem[612] = 16'h6c08;
initial mem[613] = 16'h6fe9;
initial mem[614] = 16'h7289;
initial mem[615] = 16'h746f;
initial mem[616] = 16'h75dc;
initial mem[617] = 16'h76fa;
initial mem[618] = 16'h77df;
initial mem[619] = 16'h789b;
initial mem[620] = 16'h7938;
initial mem[621] = 16'h79bd;
initial mem[622] = 16'h7a2f;
initial mem[623] = 16'h7a92;
initial mem[624] = 16'h8518;
initial mem[625] = 16'h856e;
initial mem[626] = 16'h85d1;
initial mem[627] = 16'h8643;
initial mem[628] = 16'h86c8;
initial mem[629] = 16'h8765;
initial mem[630] = 16'h8821;
initial mem[631] = 16'h8906;
initial mem[632] = 16'h8a24;
initial mem[633] = 16'h8b91;
initial mem[634] = 16'h8d77;
initial mem[635] = 16'h9017;
initial mem[636] = 16'h93f8;
initial mem[637] = 16'h9a39;
initial mem[638] = 16'ha5c9;
initial mem[639] = 16'hc001;
initial mem[640] = 16'h0;
initial mem[641] = 16'h7fff;
initial mem[642] = 16'h7fff;
initial mem[643] = 16'h7fff;
initial mem[644] = 16'h7fff;
initial mem[645] = 16'h7fff;
initial mem[646] = 16'h7fff;
initial mem[647] = 16'h7fff;
initial mem[648] = 16'h7fff;
initial mem[649] = 16'h7fff;
initial mem[650] = 16'h7fff;
initial mem[651] = 16'h7fff;
initial mem[652] = 16'h7fff;
initial mem[653] = 16'h7fff;
initial mem[654] = 16'h7fff;
initial mem[655] = 16'h7fff;
initial mem[656] = 16'h8001;
initial mem[657] = 16'h8001;
initial mem[658] = 16'h8001;
initial mem[659] = 16'h8001;
initial mem[660] = 16'h8001;
initial mem[661] = 16'h8001;
initial mem[662] = 16'h8001;
initial mem[663] = 16'h8001;
initial mem[664] = 16'h8001;
initial mem[665] = 16'h8001;
initial mem[666] = 16'h8001;
initial mem[667] = 16'h8001;
initial mem[668] = 16'h8001;
initial mem[669] = 16'h8001;
initial mem[670] = 16'h8001;
initial mem[671] = 16'h8001;
initial mem[672] = 16'h0;
initial mem[673] = 16'h3fff;
initial mem[674] = 16'h5a37;
initial mem[675] = 16'h65c7;
initial mem[676] = 16'h6c08;
initial mem[677] = 16'h6fe9;
initial mem[678] = 16'h7289;
initial mem[679] = 16'h746f;
initial mem[680] = 16'h75dc;
initial mem[681] = 16'h76fa;
initial mem[682] = 16'h77df;
initial mem[683] = 16'h789b;
initial mem[684] = 16'h7938;
initial mem[685] = 16'h79bd;
initial mem[686] = 16'h7a2f;
initial mem[687] = 16'h7a92;
initial mem[688] = 16'h8518;
initial mem[689] = 16'h856e;
initial mem[690] = 16'h85d1;
initial mem[691] = 16'h8643;
initial mem[692] = 16'h86c8;
initial mem[693] = 16'h8765;
initial mem[694] = 16'h8821;
initial mem[695] = 16'h8906;
initial mem[696] = 16'h8a24;
initial mem[697] = 16'h8b91;
initial mem[698] = 16'h8d77;
initial mem[699] = 16'h9017;
initial mem[700] = 16'h93f8;
initial mem[701] = 16'h9a39;
initial mem[702] = 16'ha5c9;
initial mem[703] = 16'hc001;
initial mem[704] = 16'h0;
initial mem[705] = 16'h7fff;
initial mem[706] = 16'h7fff;
initial mem[707] = 16'h7fff;
initial mem[708] = 16'h7fff;
initial mem[709] = 16'h7fff;
initial mem[710] = 16'h7fff;
initial mem[711] = 16'h7fff;
initial mem[712] = 16'h7fff;
initial mem[713] = 16'h7fff;
initial mem[714] = 16'h7fff;
initial mem[715] = 16'h7fff;
initial mem[716] = 16'h7fff;
initial mem[717] = 16'h7fff;
initial mem[718] = 16'h7fff;
initial mem[719] = 16'h7fff;
initial mem[720] = 16'h8001;
initial mem[721] = 16'h8001;
initial mem[722] = 16'h8001;
initial mem[723] = 16'h8001;
initial mem[724] = 16'h8001;
initial mem[725] = 16'h8001;
initial mem[726] = 16'h8001;
initial mem[727] = 16'h8001;
initial mem[728] = 16'h8001;
initial mem[729] = 16'h8001;
initial mem[730] = 16'h8001;
initial mem[731] = 16'h8001;
initial mem[732] = 16'h8001;
initial mem[733] = 16'h8001;
initial mem[734] = 16'h8001;
initial mem[735] = 16'h8001;
initial mem[736] = 16'h0;
initial mem[737] = 16'h3fff;
initial mem[738] = 16'h5a37;
initial mem[739] = 16'h65c7;
initial mem[740] = 16'h6c08;
initial mem[741] = 16'h6fe9;
initial mem[742] = 16'h7289;
initial mem[743] = 16'h746f;
initial mem[744] = 16'h75dc;
initial mem[745] = 16'h76fa;
initial mem[746] = 16'h77df;
initial mem[747] = 16'h789b;
initial mem[748] = 16'h7938;
initial mem[749] = 16'h79bd;
initial mem[750] = 16'h7a2f;
initial mem[751] = 16'h7a92;
initial mem[752] = 16'h8518;
initial mem[753] = 16'h856e;
initial mem[754] = 16'h85d1;
initial mem[755] = 16'h8643;
initial mem[756] = 16'h86c8;
initial mem[757] = 16'h8765;
initial mem[758] = 16'h8821;
initial mem[759] = 16'h8906;
initial mem[760] = 16'h8a24;
initial mem[761] = 16'h8b91;
initial mem[762] = 16'h8d77;
initial mem[763] = 16'h9017;
initial mem[764] = 16'h93f8;
initial mem[765] = 16'h9a39;
initial mem[766] = 16'ha5c9;
initial mem[767] = 16'hc001;
initial mem[768] = 16'h0;
initial mem[769] = 16'h7fff;
initial mem[770] = 16'h7fff;
initial mem[771] = 16'h7fff;
initial mem[772] = 16'h7fff;
initial mem[773] = 16'h7fff;
initial mem[774] = 16'h7fff;
initial mem[775] = 16'h7fff;
initial mem[776] = 16'h7fff;
initial mem[777] = 16'h7fff;
initial mem[778] = 16'h7fff;
initial mem[779] = 16'h7fff;
initial mem[780] = 16'h7fff;
initial mem[781] = 16'h7fff;
initial mem[782] = 16'h7fff;
initial mem[783] = 16'h7fff;
initial mem[784] = 16'h8001;
initial mem[785] = 16'h8001;
initial mem[786] = 16'h8001;
initial mem[787] = 16'h8001;
initial mem[788] = 16'h8001;
initial mem[789] = 16'h8001;
initial mem[790] = 16'h8001;
initial mem[791] = 16'h8001;
initial mem[792] = 16'h8001;
initial mem[793] = 16'h8001;
initial mem[794] = 16'h8001;
initial mem[795] = 16'h8001;
initial mem[796] = 16'h8001;
initial mem[797] = 16'h8001;
initial mem[798] = 16'h8001;
initial mem[799] = 16'h8001;
initial mem[800] = 16'h0;
initial mem[801] = 16'h3fff;
initial mem[802] = 16'h5a37;
initial mem[803] = 16'h65c7;
initial mem[804] = 16'h6c08;
initial mem[805] = 16'h6fe9;
initial mem[806] = 16'h7289;
initial mem[807] = 16'h746f;
initial mem[808] = 16'h75dc;
initial mem[809] = 16'h76fa;
initial mem[810] = 16'h77df;
initial mem[811] = 16'h789b;
initial mem[812] = 16'h7938;
initial mem[813] = 16'h79bd;
initial mem[814] = 16'h7a2f;
initial mem[815] = 16'h7a92;
initial mem[816] = 16'h8518;
initial mem[817] = 16'h856e;
initial mem[818] = 16'h85d1;
initial mem[819] = 16'h8643;
initial mem[820] = 16'h86c8;
initial mem[821] = 16'h8765;
initial mem[822] = 16'h8821;
initial mem[823] = 16'h8906;
initial mem[824] = 16'h8a24;
initial mem[825] = 16'h8b91;
initial mem[826] = 16'h8d77;
initial mem[827] = 16'h9017;
initial mem[828] = 16'h93f8;
initial mem[829] = 16'h9a39;
initial mem[830] = 16'ha5c9;
initial mem[831] = 16'hc001;
initial mem[832] = 16'h0;
initial mem[833] = 16'h7fff;
initial mem[834] = 16'h7fff;
initial mem[835] = 16'h7fff;
initial mem[836] = 16'h7fff;
initial mem[837] = 16'h7fff;
initial mem[838] = 16'h7fff;
initial mem[839] = 16'h7fff;
initial mem[840] = 16'h7fff;
initial mem[841] = 16'h7fff;
initial mem[842] = 16'h7fff;
initial mem[843] = 16'h7fff;
initial mem[844] = 16'h7fff;
initial mem[845] = 16'h7fff;
initial mem[846] = 16'h7fff;
initial mem[847] = 16'h7fff;
initial mem[848] = 16'h8001;
initial mem[849] = 16'h8001;
initial mem[850] = 16'h8001;
initial mem[851] = 16'h8001;
initial mem[852] = 16'h8001;
initial mem[853] = 16'h8001;
initial mem[854] = 16'h8001;
initial mem[855] = 16'h8001;
initial mem[856] = 16'h8001;
initial mem[857] = 16'h8001;
initial mem[858] = 16'h8001;
initial mem[859] = 16'h8001;
initial mem[860] = 16'h8001;
initial mem[861] = 16'h8001;
initial mem[862] = 16'h8001;
initial mem[863] = 16'h8001;
initial mem[864] = 16'h0;
initial mem[865] = 16'h3fff;
initial mem[866] = 16'h5a37;
initial mem[867] = 16'h65c7;
initial mem[868] = 16'h6c08;
initial mem[869] = 16'h6fe9;
initial mem[870] = 16'h7289;
initial mem[871] = 16'h746f;
initial mem[872] = 16'h75dc;
initial mem[873] = 16'h76fa;
initial mem[874] = 16'h77df;
initial mem[875] = 16'h789b;
initial mem[876] = 16'h7938;
initial mem[877] = 16'h79bd;
initial mem[878] = 16'h7a2f;
initial mem[879] = 16'h7a92;
initial mem[880] = 16'h8518;
initial mem[881] = 16'h856e;
initial mem[882] = 16'h85d1;
initial mem[883] = 16'h8643;
initial mem[884] = 16'h86c8;
initial mem[885] = 16'h8765;
initial mem[886] = 16'h8821;
initial mem[887] = 16'h8906;
initial mem[888] = 16'h8a24;
initial mem[889] = 16'h8b91;
initial mem[890] = 16'h8d77;
initial mem[891] = 16'h9017;
initial mem[892] = 16'h93f8;
initial mem[893] = 16'h9a39;
initial mem[894] = 16'ha5c9;
initial mem[895] = 16'hc001;
initial mem[896] = 16'h0;
initial mem[897] = 16'h7fff;
initial mem[898] = 16'h7fff;
initial mem[899] = 16'h7fff;
initial mem[900] = 16'h7fff;
initial mem[901] = 16'h7fff;
initial mem[902] = 16'h7fff;
initial mem[903] = 16'h7fff;
initial mem[904] = 16'h7fff;
initial mem[905] = 16'h7fff;
initial mem[906] = 16'h7fff;
initial mem[907] = 16'h7fff;
initial mem[908] = 16'h7fff;
initial mem[909] = 16'h7fff;
initial mem[910] = 16'h7fff;
initial mem[911] = 16'h7fff;
initial mem[912] = 16'h8001;
initial mem[913] = 16'h8001;
initial mem[914] = 16'h8001;
initial mem[915] = 16'h8001;
initial mem[916] = 16'h8001;
initial mem[917] = 16'h8001;
initial mem[918] = 16'h8001;
initial mem[919] = 16'h8001;
initial mem[920] = 16'h8001;
initial mem[921] = 16'h8001;
initial mem[922] = 16'h8001;
initial mem[923] = 16'h8001;
initial mem[924] = 16'h8001;
initial mem[925] = 16'h8001;
initial mem[926] = 16'h8001;
initial mem[927] = 16'h8001;
initial mem[928] = 16'h0;
initial mem[929] = 16'h3fff;
initial mem[930] = 16'h5a37;
initial mem[931] = 16'h65c7;
initial mem[932] = 16'h6c08;
initial mem[933] = 16'h6fe9;
initial mem[934] = 16'h7289;
initial mem[935] = 16'h746f;
initial mem[936] = 16'h75dc;
initial mem[937] = 16'h76fa;
initial mem[938] = 16'h77df;
initial mem[939] = 16'h789b;
initial mem[940] = 16'h7938;
initial mem[941] = 16'h79bd;
initial mem[942] = 16'h7a2f;
initial mem[943] = 16'h7a92;
initial mem[944] = 16'h8518;
initial mem[945] = 16'h856e;
initial mem[946] = 16'h85d1;
initial mem[947] = 16'h8643;
initial mem[948] = 16'h86c8;
initial mem[949] = 16'h8765;
initial mem[950] = 16'h8821;
initial mem[951] = 16'h8906;
initial mem[952] = 16'h8a24;
initial mem[953] = 16'h8b91;
initial mem[954] = 16'h8d77;
initial mem[955] = 16'h9017;
initial mem[956] = 16'h93f8;
initial mem[957] = 16'h9a39;
initial mem[958] = 16'ha5c9;
initial mem[959] = 16'hc001;
initial mem[960] = 16'h0;
initial mem[961] = 16'h7fff;
initial mem[962] = 16'h7fff;
initial mem[963] = 16'h7fff;
initial mem[964] = 16'h7fff;
initial mem[965] = 16'h7fff;
initial mem[966] = 16'h7fff;
initial mem[967] = 16'h7fff;
initial mem[968] = 16'h7fff;
initial mem[969] = 16'h7fff;
initial mem[970] = 16'h7fff;
initial mem[971] = 16'h7fff;
initial mem[972] = 16'h7fff;
initial mem[973] = 16'h7fff;
initial mem[974] = 16'h7fff;
initial mem[975] = 16'h7fff;
initial mem[976] = 16'h8001;
initial mem[977] = 16'h8001;
initial mem[978] = 16'h8001;
initial mem[979] = 16'h8001;
initial mem[980] = 16'h8001;
initial mem[981] = 16'h8001;
initial mem[982] = 16'h8001;
initial mem[983] = 16'h8001;
initial mem[984] = 16'h8001;
initial mem[985] = 16'h8001;
initial mem[986] = 16'h8001;
initial mem[987] = 16'h8001;
initial mem[988] = 16'h8001;
initial mem[989] = 16'h8001;
initial mem[990] = 16'h8001;
initial mem[991] = 16'h8001;
initial mem[992] = 16'h0;
initial mem[993] = 16'h3fff;
initial mem[994] = 16'h5a37;
initial mem[995] = 16'h65c7;
initial mem[996] = 16'h6c08;
initial mem[997] = 16'h6fe9;
initial mem[998] = 16'h7289;
initial mem[999] = 16'h746f;
initial mem[1000] = 16'h75dc;
initial mem[1001] = 16'h76fa;
initial mem[1002] = 16'h77df;
initial mem[1003] = 16'h789b;
initial mem[1004] = 16'h7938;
initial mem[1005] = 16'h79bd;
initial mem[1006] = 16'h7a2f;
initial mem[1007] = 16'h7a92;
initial mem[1008] = 16'h8518;
initial mem[1009] = 16'h856e;
initial mem[1010] = 16'h85d1;
initial mem[1011] = 16'h8643;
initial mem[1012] = 16'h86c8;
initial mem[1013] = 16'h8765;
initial mem[1014] = 16'h8821;
initial mem[1015] = 16'h8906;
initial mem[1016] = 16'h8a24;
initial mem[1017] = 16'h8b91;
initial mem[1018] = 16'h8d77;
initial mem[1019] = 16'h9017;
initial mem[1020] = 16'h93f8;
initial mem[1021] = 16'h9a39;
initial mem[1022] = 16'ha5c9;
initial mem[1023] = 16'hc001;
always @(posedge clk) begin
	data <= mem[addr];
end
endmodule
