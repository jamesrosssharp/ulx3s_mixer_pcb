module vuTable(input clk, input [9:0] addr, output reg [7:0] data);
reg [15:0] mem [0:1023];
initial mem[0] = 8'h0;
initial mem[1] = 8'h0;
initial mem[2] = 8'h0;
initial mem[3] = 8'h0;
initial mem[4] = 8'h0;
initial mem[5] = 8'h0;
initial mem[6] = 8'h0;
initial mem[7] = 8'h0;
initial mem[8] = 8'h0;
initial mem[9] = 8'h0;
initial mem[10] = 8'h0;
initial mem[11] = 8'h0;
initial mem[12] = 8'h0;
initial mem[13] = 8'h0;
initial mem[14] = 8'h0;
initial mem[15] = 8'h0;
initial mem[16] = 8'h0;
initial mem[17] = 8'h0;
initial mem[18] = 8'h0;
initial mem[19] = 8'h0;
initial mem[20] = 8'h0;
initial mem[21] = 8'h0;
initial mem[22] = 8'h0;
initial mem[23] = 8'h0;
initial mem[24] = 8'h0;
initial mem[25] = 8'h0;
initial mem[26] = 8'h0;
initial mem[27] = 8'h0;
initial mem[28] = 8'h0;
initial mem[29] = 8'h0;
initial mem[30] = 8'h0;
initial mem[31] = 8'h0;
initial mem[32] = 8'h0;
initial mem[33] = 8'h0;
initial mem[34] = 8'h0;
initial mem[35] = 8'h0;
initial mem[36] = 8'h0;
initial mem[37] = 8'h0;
initial mem[38] = 8'h0;
initial mem[39] = 8'h0;
initial mem[40] = 8'h0;
initial mem[41] = 8'h0;
initial mem[42] = 8'h0;
initial mem[43] = 8'h0;
initial mem[44] = 8'h0;
initial mem[45] = 8'h0;
initial mem[46] = 8'h0;
initial mem[47] = 8'h0;
initial mem[48] = 8'h0;
initial mem[49] = 8'h0;
initial mem[50] = 8'h0;
initial mem[51] = 8'h0;
initial mem[52] = 8'h0;
initial mem[53] = 8'h0;
initial mem[54] = 8'h0;
initial mem[55] = 8'h0;
initial mem[56] = 8'h0;
initial mem[57] = 8'h0;
initial mem[58] = 8'h0;
initial mem[59] = 8'h0;
initial mem[60] = 8'h0;
initial mem[61] = 8'h0;
initial mem[62] = 8'h0;
initial mem[63] = 8'h0;
initial mem[64] = 8'h0;
initial mem[65] = 8'h0;
initial mem[66] = 8'h0;
initial mem[67] = 8'h0;
initial mem[68] = 8'h0;
initial mem[69] = 8'h0;
initial mem[70] = 8'h0;
initial mem[71] = 8'h0;
initial mem[72] = 8'h0;
initial mem[73] = 8'h0;
initial mem[74] = 8'h0;
initial mem[75] = 8'h0;
initial mem[76] = 8'h0;
initial mem[77] = 8'h0;
initial mem[78] = 8'h0;
initial mem[79] = 8'h0;
initial mem[80] = 8'h0;
initial mem[81] = 8'h0;
initial mem[82] = 8'h0;
initial mem[83] = 8'h0;
initial mem[84] = 8'h0;
initial mem[85] = 8'h0;
initial mem[86] = 8'h0;
initial mem[87] = 8'h0;
initial mem[88] = 8'h0;
initial mem[89] = 8'h0;
initial mem[90] = 8'h0;
initial mem[91] = 8'h0;
initial mem[92] = 8'h0;
initial mem[93] = 8'h0;
initial mem[94] = 8'h0;
initial mem[95] = 8'h0;
initial mem[96] = 8'h0;
initial mem[97] = 8'h0;
initial mem[98] = 8'h0;
initial mem[99] = 8'h0;
initial mem[100] = 8'h0;
initial mem[101] = 8'h0;
initial mem[102] = 8'h0;
initial mem[103] = 8'h0;
initial mem[104] = 8'h0;
initial mem[105] = 8'h0;
initial mem[106] = 8'h0;
initial mem[107] = 8'h0;
initial mem[108] = 8'h0;
initial mem[109] = 8'h0;
initial mem[110] = 8'h0;
initial mem[111] = 8'h0;
initial mem[112] = 8'h0;
initial mem[113] = 8'h0;
initial mem[114] = 8'h0;
initial mem[115] = 8'h0;
initial mem[116] = 8'h0;
initial mem[117] = 8'h0;
initial mem[118] = 8'h0;
initial mem[119] = 8'h0;
initial mem[120] = 8'h1;
initial mem[121] = 8'h1;
initial mem[122] = 8'h1;
initial mem[123] = 8'h1;
initial mem[124] = 8'h1;
initial mem[125] = 8'h1;
initial mem[126] = 8'h1;
initial mem[127] = 8'h1;
initial mem[128] = 8'h1;
initial mem[129] = 8'h1;
initial mem[130] = 8'h1;
initial mem[131] = 8'h1;
initial mem[132] = 8'h1;
initial mem[133] = 8'h1;
initial mem[134] = 8'h1;
initial mem[135] = 8'h1;
initial mem[136] = 8'h1;
initial mem[137] = 8'h1;
initial mem[138] = 8'h1;
initial mem[139] = 8'h1;
initial mem[140] = 8'h1;
initial mem[141] = 8'h1;
initial mem[142] = 8'h1;
initial mem[143] = 8'h1;
initial mem[144] = 8'h1;
initial mem[145] = 8'h1;
initial mem[146] = 8'h1;
initial mem[147] = 8'h1;
initial mem[148] = 8'h1;
initial mem[149] = 8'h1;
initial mem[150] = 8'h1;
initial mem[151] = 8'h1;
initial mem[152] = 8'h1;
initial mem[153] = 8'h1;
initial mem[154] = 8'h1;
initial mem[155] = 8'h1;
initial mem[156] = 8'h1;
initial mem[157] = 8'h1;
initial mem[158] = 8'h1;
initial mem[159] = 8'h1;
initial mem[160] = 8'h1;
initial mem[161] = 8'h1;
initial mem[162] = 8'h1;
initial mem[163] = 8'h1;
initial mem[164] = 8'h1;
initial mem[165] = 8'h1;
initial mem[166] = 8'h1;
initial mem[167] = 8'h1;
initial mem[168] = 8'h1;
initial mem[169] = 8'h1;
initial mem[170] = 8'h1;
initial mem[171] = 8'h1;
initial mem[172] = 8'h1;
initial mem[173] = 8'h1;
initial mem[174] = 8'h1;
initial mem[175] = 8'h1;
initial mem[176] = 8'h1;
initial mem[177] = 8'h1;
initial mem[178] = 8'h1;
initial mem[179] = 8'h1;
initial mem[180] = 8'h1;
initial mem[181] = 8'h1;
initial mem[182] = 8'h1;
initial mem[183] = 8'h1;
initial mem[184] = 8'h1;
initial mem[185] = 8'h1;
initial mem[186] = 8'h1;
initial mem[187] = 8'h1;
initial mem[188] = 8'h1;
initial mem[189] = 8'h1;
initial mem[190] = 8'h1;
initial mem[191] = 8'h1;
initial mem[192] = 8'h1;
initial mem[193] = 8'h1;
initial mem[194] = 8'h1;
initial mem[195] = 8'h1;
initial mem[196] = 8'h1;
initial mem[197] = 8'h1;
initial mem[198] = 8'h1;
initial mem[199] = 8'h1;
initial mem[200] = 8'hf;
initial mem[201] = 8'hf;
initial mem[202] = 8'hf;
initial mem[203] = 8'hf;
initial mem[204] = 8'hf;
initial mem[205] = 8'hf;
initial mem[206] = 8'hf;
initial mem[207] = 8'hf;
initial mem[208] = 8'hf;
initial mem[209] = 8'hf;
initial mem[210] = 8'hf;
initial mem[211] = 8'hf;
initial mem[212] = 8'hf;
initial mem[213] = 8'hf;
initial mem[214] = 8'hf;
initial mem[215] = 8'hf;
initial mem[216] = 8'hf;
initial mem[217] = 8'hf;
initial mem[218] = 8'hf;
initial mem[219] = 8'hf;
initial mem[220] = 8'hf;
initial mem[221] = 8'hf;
initial mem[222] = 8'hf;
initial mem[223] = 8'hf;
initial mem[224] = 8'hf;
initial mem[225] = 8'hf;
initial mem[226] = 8'hf;
initial mem[227] = 8'hf;
initial mem[228] = 8'hf;
initial mem[229] = 8'hf;
initial mem[230] = 8'hf;
initial mem[231] = 8'hf;
initial mem[232] = 8'hf;
initial mem[233] = 8'hf;
initial mem[234] = 8'hf;
initial mem[235] = 8'hf;
initial mem[236] = 8'hf;
initial mem[237] = 8'hf;
initial mem[238] = 8'hf;
initial mem[239] = 8'hf;
initial mem[240] = 8'hf;
initial mem[241] = 8'hf;
initial mem[242] = 8'hf;
initial mem[243] = 8'hf;
initial mem[244] = 8'hf;
initial mem[245] = 8'hf;
initial mem[246] = 8'hf;
initial mem[247] = 8'hf;
initial mem[248] = 8'hf;
initial mem[249] = 8'hf;
initial mem[250] = 8'hf;
initial mem[251] = 8'hf;
initial mem[252] = 8'hf;
initial mem[253] = 8'hf;
initial mem[254] = 8'hf;
initial mem[255] = 8'hf;
initial mem[256] = 8'hf;
initial mem[257] = 8'hf;
initial mem[258] = 8'hf;
initial mem[259] = 8'hf;
initial mem[260] = 8'hf;
initial mem[261] = 8'hf;
initial mem[262] = 8'hf;
initial mem[263] = 8'hf;
initial mem[264] = 8'hf;
initial mem[265] = 8'hf;
initial mem[266] = 8'hf;
initial mem[267] = 8'hf;
initial mem[268] = 8'hf;
initial mem[269] = 8'hf;
initial mem[270] = 8'hf;
initial mem[271] = 8'hf;
initial mem[272] = 8'hf;
initial mem[273] = 8'hf;
initial mem[274] = 8'hf;
initial mem[275] = 8'hf;
initial mem[276] = 8'hf;
initial mem[277] = 8'hf;
initial mem[278] = 8'hf;
initial mem[279] = 8'hf;
initial mem[280] = 8'hf;
initial mem[281] = 8'hf;
initial mem[282] = 8'hf;
initial mem[283] = 8'hf;
initial mem[284] = 8'hf;
initial mem[285] = 8'hf;
initial mem[286] = 8'hf;
initial mem[287] = 8'hf;
initial mem[288] = 8'hf;
initial mem[289] = 8'hf;
initial mem[290] = 8'hf;
initial mem[291] = 8'hf;
initial mem[292] = 8'hf;
initial mem[293] = 8'hf;
initial mem[294] = 8'hf;
initial mem[295] = 8'hf;
initial mem[296] = 8'hf;
initial mem[297] = 8'hf;
initial mem[298] = 8'hf;
initial mem[299] = 8'hf;
initial mem[300] = 8'hf;
initial mem[301] = 8'hf;
initial mem[302] = 8'hf;
initial mem[303] = 8'hf;
initial mem[304] = 8'hf;
initial mem[305] = 8'hf;
initial mem[306] = 8'hf;
initial mem[307] = 8'hf;
initial mem[308] = 8'hf;
initial mem[309] = 8'hf;
initial mem[310] = 8'hf;
initial mem[311] = 8'hf;
initial mem[312] = 8'hf;
initial mem[313] = 8'hf;
initial mem[314] = 8'hf;
initial mem[315] = 8'hf;
initial mem[316] = 8'hf;
initial mem[317] = 8'hf;
initial mem[318] = 8'hf;
initial mem[319] = 8'hf;
initial mem[320] = 8'hf;
initial mem[321] = 8'hf;
initial mem[322] = 8'hf;
initial mem[323] = 8'hf;
initial mem[324] = 8'hf;
initial mem[325] = 8'hf;
initial mem[326] = 8'hf;
initial mem[327] = 8'hf;
initial mem[328] = 8'hf;
initial mem[329] = 8'hf;
initial mem[330] = 8'hf;
initial mem[331] = 8'hf;
initial mem[332] = 8'hf;
initial mem[333] = 8'hf;
initial mem[334] = 8'hf;
initial mem[335] = 8'hf;
initial mem[336] = 8'hf;
initial mem[337] = 8'hf;
initial mem[338] = 8'hf;
initial mem[339] = 8'hf;
initial mem[340] = 8'hf;
initial mem[341] = 8'hf;
initial mem[342] = 8'hf;
initial mem[343] = 8'hf;
initial mem[344] = 8'hf;
initial mem[345] = 8'hf;
initial mem[346] = 8'hf;
initial mem[347] = 8'hf;
initial mem[348] = 8'hf;
initial mem[349] = 8'hf;
initial mem[350] = 8'hf;
initial mem[351] = 8'hf;
initial mem[352] = 8'hf;
initial mem[353] = 8'hf;
initial mem[354] = 8'hf;
initial mem[355] = 8'hf;
initial mem[356] = 8'hf;
initial mem[357] = 8'hf;
initial mem[358] = 8'hf;
initial mem[359] = 8'hf;
initial mem[360] = 8'hf;
initial mem[361] = 8'hf;
initial mem[362] = 8'hf;
initial mem[363] = 8'hf;
initial mem[364] = 8'hf;
initial mem[365] = 8'hf;
initial mem[366] = 8'hf;
initial mem[367] = 8'hf;
initial mem[368] = 8'hf;
initial mem[369] = 8'hf;
initial mem[370] = 8'hf;
initial mem[371] = 8'hf;
initial mem[372] = 8'hf;
initial mem[373] = 8'hf;
initial mem[374] = 8'hf;
initial mem[375] = 8'hf;
initial mem[376] = 8'hf;
initial mem[377] = 8'hf;
initial mem[378] = 8'hf;
initial mem[379] = 8'hf;
initial mem[380] = 8'hf;
initial mem[381] = 8'hf;
initial mem[382] = 8'hf;
initial mem[383] = 8'hf;
initial mem[384] = 8'hf;
initial mem[385] = 8'hf;
initial mem[386] = 8'hf;
initial mem[387] = 8'hf;
initial mem[388] = 8'hf;
initial mem[389] = 8'hf;
initial mem[390] = 8'hf;
initial mem[391] = 8'hf;
initial mem[392] = 8'hf;
initial mem[393] = 8'hf;
initial mem[394] = 8'hf;
initial mem[395] = 8'hf;
initial mem[396] = 8'hf;
initial mem[397] = 8'hf;
initial mem[398] = 8'hf;
initial mem[399] = 8'hf;
initial mem[400] = 8'hf;
initial mem[401] = 8'h3;
initial mem[402] = 8'h3;
initial mem[403] = 8'h3;
initial mem[404] = 8'h3;
initial mem[405] = 8'h3;
initial mem[406] = 8'h3;
initial mem[407] = 8'h3;
initial mem[408] = 8'h3;
initial mem[409] = 8'h3;
initial mem[410] = 8'h3;
initial mem[411] = 8'h3;
initial mem[412] = 8'h3;
initial mem[413] = 8'h3;
initial mem[414] = 8'h3;
initial mem[415] = 8'h3;
initial mem[416] = 8'h3;
initial mem[417] = 8'h3;
initial mem[418] = 8'h3;
initial mem[419] = 8'h3;
initial mem[420] = 8'h3;
initial mem[421] = 8'h3;
initial mem[422] = 8'h3;
initial mem[423] = 8'h3;
initial mem[424] = 8'h3;
initial mem[425] = 8'h3;
initial mem[426] = 8'h3;
initial mem[427] = 8'h3;
initial mem[428] = 8'h3;
initial mem[429] = 8'h3;
initial mem[430] = 8'h3;
initial mem[431] = 8'h3;
initial mem[432] = 8'h3;
initial mem[433] = 8'h3;
initial mem[434] = 8'h3;
initial mem[435] = 8'h3;
initial mem[436] = 8'h3;
initial mem[437] = 8'h3;
initial mem[438] = 8'h3;
initial mem[439] = 8'h3;
initial mem[440] = 8'h3;
initial mem[441] = 8'h3;
initial mem[442] = 8'h3;
initial mem[443] = 8'h3;
initial mem[444] = 8'h3;
initial mem[445] = 8'h3;
initial mem[446] = 8'h3;
initial mem[447] = 8'h3;
initial mem[448] = 8'h3;
initial mem[449] = 8'h3;
initial mem[450] = 8'h3;
initial mem[451] = 8'h3;
initial mem[452] = 8'h3;
initial mem[453] = 8'h3;
initial mem[454] = 8'h3;
initial mem[455] = 8'h3;
initial mem[456] = 8'h3;
initial mem[457] = 8'h3;
initial mem[458] = 8'h3;
initial mem[459] = 8'h3;
initial mem[460] = 8'h3;
initial mem[461] = 8'h3;
initial mem[462] = 8'h3;
initial mem[463] = 8'h3;
initial mem[464] = 8'h3;
initial mem[465] = 8'h3;
initial mem[466] = 8'h3;
initial mem[467] = 8'h3;
initial mem[468] = 8'h3;
initial mem[469] = 8'h3;
initial mem[470] = 8'h3;
initial mem[471] = 8'h3;
initial mem[472] = 8'h3;
initial mem[473] = 8'h3;
initial mem[474] = 8'h3;
initial mem[475] = 8'h3;
initial mem[476] = 8'h3;
initial mem[477] = 8'h3;
initial mem[478] = 8'h3;
initial mem[479] = 8'h3;
initial mem[480] = 8'h3;
initial mem[481] = 8'h3;
initial mem[482] = 8'h3;
initial mem[483] = 8'h3;
initial mem[484] = 8'h3;
initial mem[485] = 8'h3;
initial mem[486] = 8'h3;
initial mem[487] = 8'h3;
initial mem[488] = 8'h3;
initial mem[489] = 8'h3;
initial mem[490] = 8'h3;
initial mem[491] = 8'h3;
initial mem[492] = 8'h3;
initial mem[493] = 8'h3;
initial mem[494] = 8'h3;
initial mem[495] = 8'h3;
initial mem[496] = 8'h3;
initial mem[497] = 8'h3;
initial mem[498] = 8'h3;
initial mem[499] = 8'h3;
initial mem[500] = 8'h3;
initial mem[501] = 8'h3;
initial mem[502] = 8'h3;
initial mem[503] = 8'h3;
initial mem[504] = 8'h3;
initial mem[505] = 8'h3;
initial mem[506] = 8'h3;
initial mem[507] = 8'h3;
initial mem[508] = 8'h3;
initial mem[509] = 8'h3;
initial mem[510] = 8'h3;
initial mem[511] = 8'h3;
initial mem[512] = 8'h3;
initial mem[513] = 8'h3;
initial mem[514] = 8'h3;
initial mem[515] = 8'h3;
initial mem[516] = 8'h3;
initial mem[517] = 8'h3;
initial mem[518] = 8'h3;
initial mem[519] = 8'h3;
initial mem[520] = 8'h3;
initial mem[521] = 8'h3;
initial mem[522] = 8'h3;
initial mem[523] = 8'h3;
initial mem[524] = 8'h3;
initial mem[525] = 8'h3;
initial mem[526] = 8'h3;
initial mem[527] = 8'h3;
initial mem[528] = 8'h3;
initial mem[529] = 8'h3;
initial mem[530] = 8'h3;
initial mem[531] = 8'h3;
initial mem[532] = 8'h3;
initial mem[533] = 8'h3;
initial mem[534] = 8'h3;
initial mem[535] = 8'h3;
initial mem[536] = 8'h3;
initial mem[537] = 8'h3;
initial mem[538] = 8'h3;
initial mem[539] = 8'h3;
initial mem[540] = 8'h3;
initial mem[541] = 8'h3;
initial mem[542] = 8'h3;
initial mem[543] = 8'h3;
initial mem[544] = 8'h3;
initial mem[545] = 8'h3;
initial mem[546] = 8'h3;
initial mem[547] = 8'h3;
initial mem[548] = 8'h3;
initial mem[549] = 8'h3;
initial mem[550] = 8'h3;
initial mem[551] = 8'h3;
initial mem[552] = 8'h3;
initial mem[553] = 8'h3;
initial mem[554] = 8'h3;
initial mem[555] = 8'h3;
initial mem[556] = 8'h3;
initial mem[557] = 8'h3;
initial mem[558] = 8'h3;
initial mem[559] = 8'h3;
initial mem[560] = 8'h3;
initial mem[561] = 8'h3;
initial mem[562] = 8'h3;
initial mem[563] = 8'h3;
initial mem[564] = 8'h3;
initial mem[565] = 8'h3;
initial mem[566] = 8'h3;
initial mem[567] = 8'h3;
initial mem[568] = 8'h3;
initial mem[569] = 8'h3;
initial mem[570] = 8'h3;
initial mem[571] = 8'h3;
initial mem[572] = 8'h3;
initial mem[573] = 8'h3;
initial mem[574] = 8'h3;
initial mem[575] = 8'h3;
initial mem[576] = 8'h3;
initial mem[577] = 8'h3;
initial mem[578] = 8'h3;
initial mem[579] = 8'h3;
initial mem[580] = 8'h3;
initial mem[581] = 8'h3;
initial mem[582] = 8'h3;
initial mem[583] = 8'h3;
initial mem[584] = 8'h3;
initial mem[585] = 8'h3;
initial mem[586] = 8'h3;
initial mem[587] = 8'h3;
initial mem[588] = 8'h3;
initial mem[589] = 8'h3;
initial mem[590] = 8'h3;
initial mem[591] = 8'h3;
initial mem[592] = 8'h3;
initial mem[593] = 8'h3;
initial mem[594] = 8'h3;
initial mem[595] = 8'h3;
initial mem[596] = 8'h3;
initial mem[597] = 8'h3;
initial mem[598] = 8'h3;
initial mem[599] = 8'h3;
initial mem[600] = 8'h3;
initial mem[601] = 8'h3;
initial mem[602] = 8'h3;
initial mem[603] = 8'h3;
initial mem[604] = 8'h3;
initial mem[605] = 8'h3;
initial mem[606] = 8'h3;
initial mem[607] = 8'h3;
initial mem[608] = 8'h3;
initial mem[609] = 8'h3;
initial mem[610] = 8'h3;
initial mem[611] = 8'h3;
initial mem[612] = 8'h3;
initial mem[613] = 8'h3;
initial mem[614] = 8'h3;
initial mem[615] = 8'h3;
initial mem[616] = 8'h3;
initial mem[617] = 8'h3;
initial mem[618] = 8'h3;
initial mem[619] = 8'h3;
initial mem[620] = 8'h3;
initial mem[621] = 8'h3;
initial mem[622] = 8'h3;
initial mem[623] = 8'h3;
initial mem[624] = 8'h3;
initial mem[625] = 8'h3;
initial mem[626] = 8'h3;
initial mem[627] = 8'h3;
initial mem[628] = 8'h3;
initial mem[629] = 8'h3;
initial mem[630] = 8'h3;
initial mem[631] = 8'h3;
initial mem[632] = 8'h3;
initial mem[633] = 8'h3;
initial mem[634] = 8'h3;
initial mem[635] = 8'h3;
initial mem[636] = 8'h3;
initial mem[637] = 8'h3;
initial mem[638] = 8'h3;
initial mem[639] = 8'h3;
initial mem[640] = 8'h3;
initial mem[641] = 8'h3;
initial mem[642] = 8'h3;
initial mem[643] = 8'h3;
initial mem[644] = 8'h3;
initial mem[645] = 8'h3;
initial mem[646] = 8'h3;
initial mem[647] = 8'h3;
initial mem[648] = 8'h3;
initial mem[649] = 8'h3;
initial mem[650] = 8'h3;
initial mem[651] = 8'h3;
initial mem[652] = 8'h3;
initial mem[653] = 8'h3;
initial mem[654] = 8'h3;
initial mem[655] = 8'h3;
initial mem[656] = 8'h3;
initial mem[657] = 8'h3;
initial mem[658] = 8'h3;
initial mem[659] = 8'h3;
initial mem[660] = 8'h3;
initial mem[661] = 8'h3;
initial mem[662] = 8'h3;
initial mem[663] = 8'h3;
initial mem[664] = 8'h3;
initial mem[665] = 8'h3;
initial mem[666] = 8'h3;
initial mem[667] = 8'h3;
initial mem[668] = 8'h3;
initial mem[669] = 8'h3;
initial mem[670] = 8'h3;
initial mem[671] = 8'h3;
initial mem[672] = 8'h3;
initial mem[673] = 8'h3;
initial mem[674] = 8'h3;
initial mem[675] = 8'h3;
initial mem[676] = 8'h3;
initial mem[677] = 8'h3;
initial mem[678] = 8'h3;
initial mem[679] = 8'h3;
initial mem[680] = 8'h3;
initial mem[681] = 8'h3;
initial mem[682] = 8'h3;
initial mem[683] = 8'h3;
initial mem[684] = 8'h3;
initial mem[685] = 8'h3;
initial mem[686] = 8'h3;
initial mem[687] = 8'h3;
initial mem[688] = 8'h3;
initial mem[689] = 8'h3;
initial mem[690] = 8'h3;
initial mem[691] = 8'h3;
initial mem[692] = 8'h3;
initial mem[693] = 8'h3;
initial mem[694] = 8'h3;
initial mem[695] = 8'h3;
initial mem[696] = 8'h3;
initial mem[697] = 8'h3;
initial mem[698] = 8'h3;
initial mem[699] = 8'h3;
initial mem[700] = 8'h3;
initial mem[701] = 8'h3;
initial mem[702] = 8'h3;
initial mem[703] = 8'h3;
initial mem[704] = 8'h3;
initial mem[705] = 8'h3;
initial mem[706] = 8'h3;
initial mem[707] = 8'h3;
initial mem[708] = 8'h3;
initial mem[709] = 8'h3;
initial mem[710] = 8'h3;
initial mem[711] = 8'h3;
initial mem[712] = 8'h3;
initial mem[713] = 8'h3;
initial mem[714] = 8'h3;
initial mem[715] = 8'h3;
initial mem[716] = 8'h3;
initial mem[717] = 8'h3;
initial mem[718] = 8'h3;
initial mem[719] = 8'h3;
initial mem[720] = 8'h3;
initial mem[721] = 8'h3;
initial mem[722] = 8'h3;
initial mem[723] = 8'h3;
initial mem[724] = 8'h3;
initial mem[725] = 8'h3;
initial mem[726] = 8'h3;
initial mem[727] = 8'h3;
initial mem[728] = 8'h3;
initial mem[729] = 8'h3;
initial mem[730] = 8'h3;
initial mem[731] = 8'h3;
initial mem[732] = 8'h3;
initial mem[733] = 8'h3;
initial mem[734] = 8'h3;
initial mem[735] = 8'h3;
initial mem[736] = 8'h3;
initial mem[737] = 8'h3;
initial mem[738] = 8'h3;
initial mem[739] = 8'h3;
initial mem[740] = 8'h3;
initial mem[741] = 8'h3;
initial mem[742] = 8'h3;
initial mem[743] = 8'h3;
initial mem[744] = 8'h3;
initial mem[745] = 8'h3;
initial mem[746] = 8'h3;
initial mem[747] = 8'h3;
initial mem[748] = 8'h3;
initial mem[749] = 8'h3;
initial mem[750] = 8'h3;
initial mem[751] = 8'h3;
initial mem[752] = 8'h3;
initial mem[753] = 8'h3;
initial mem[754] = 8'h3;
initial mem[755] = 8'h3;
initial mem[756] = 8'h3;
initial mem[757] = 8'h3;
initial mem[758] = 8'h3;
initial mem[759] = 8'h3;
initial mem[760] = 8'h3;
initial mem[761] = 8'h3;
initial mem[762] = 8'h3;
initial mem[763] = 8'h3;
initial mem[764] = 8'h3;
initial mem[765] = 8'h3;
initial mem[766] = 8'h3;
initial mem[767] = 8'h3;
initial mem[768] = 8'h3;
initial mem[769] = 8'h3;
initial mem[770] = 8'h3;
initial mem[771] = 8'h3;
initial mem[772] = 8'h3;
initial mem[773] = 8'h3;
initial mem[774] = 8'h3;
initial mem[775] = 8'h3;
initial mem[776] = 8'h3;
initial mem[777] = 8'h3;
initial mem[778] = 8'h3;
initial mem[779] = 8'h3;
initial mem[780] = 8'h3;
initial mem[781] = 8'h3;
initial mem[782] = 8'h3;
initial mem[783] = 8'h3;
initial mem[784] = 8'h3;
initial mem[785] = 8'h3;
initial mem[786] = 8'h3;
initial mem[787] = 8'h3;
initial mem[788] = 8'h3;
initial mem[789] = 8'h3;
initial mem[790] = 8'h3;
initial mem[791] = 8'h3;
initial mem[792] = 8'h3;
initial mem[793] = 8'h3;
initial mem[794] = 8'h3;
initial mem[795] = 8'h3;
initial mem[796] = 8'h3;
initial mem[797] = 8'h3;
initial mem[798] = 8'h3;
initial mem[799] = 8'h3;
initial mem[800] = 8'h3;
initial mem[801] = 8'h3;
initial mem[802] = 8'h3;
initial mem[803] = 8'h3;
initial mem[804] = 8'h3;
initial mem[805] = 8'h3;
initial mem[806] = 8'h3;
initial mem[807] = 8'h3;
initial mem[808] = 8'h3;
initial mem[809] = 8'h3;
initial mem[810] = 8'h3;
initial mem[811] = 8'h3;
initial mem[812] = 8'h3;
initial mem[813] = 8'h3;
initial mem[814] = 8'h3;
initial mem[815] = 8'h3;
initial mem[816] = 8'h3;
initial mem[817] = 8'h3;
initial mem[818] = 8'h3;
initial mem[819] = 8'h3;
initial mem[820] = 8'h3;
initial mem[821] = 8'h3;
initial mem[822] = 8'h3;
initial mem[823] = 8'h3;
initial mem[824] = 8'h3;
initial mem[825] = 8'h3;
initial mem[826] = 8'h3;
initial mem[827] = 8'h3;
initial mem[828] = 8'h3;
initial mem[829] = 8'h3;
initial mem[830] = 8'h3;
initial mem[831] = 8'h3;
initial mem[832] = 8'h3;
initial mem[833] = 8'h3;
initial mem[834] = 8'h3;
initial mem[835] = 8'h3;
initial mem[836] = 8'h3;
initial mem[837] = 8'h3;
initial mem[838] = 8'h3;
initial mem[839] = 8'h3;
initial mem[840] = 8'h3;
initial mem[841] = 8'h3;
initial mem[842] = 8'h3;
initial mem[843] = 8'h3;
initial mem[844] = 8'h3;
initial mem[845] = 8'h3;
initial mem[846] = 8'h3;
initial mem[847] = 8'h3;
initial mem[848] = 8'h3;
initial mem[849] = 8'h3;
initial mem[850] = 8'h3;
initial mem[851] = 8'h3;
initial mem[852] = 8'h3;
initial mem[853] = 8'h3;
initial mem[854] = 8'h3;
initial mem[855] = 8'h3;
initial mem[856] = 8'h3;
initial mem[857] = 8'h3;
initial mem[858] = 8'h3;
initial mem[859] = 8'h3;
initial mem[860] = 8'h3;
initial mem[861] = 8'h3;
initial mem[862] = 8'h3;
initial mem[863] = 8'h3;
initial mem[864] = 8'h3;
initial mem[865] = 8'h3;
initial mem[866] = 8'h3;
initial mem[867] = 8'h3;
initial mem[868] = 8'h3;
initial mem[869] = 8'h3;
initial mem[870] = 8'h3;
initial mem[871] = 8'h3;
initial mem[872] = 8'h3;
initial mem[873] = 8'h3;
initial mem[874] = 8'h3;
initial mem[875] = 8'h3;
initial mem[876] = 8'h3;
initial mem[877] = 8'h3;
initial mem[878] = 8'h3;
initial mem[879] = 8'h3;
initial mem[880] = 8'h3;
initial mem[881] = 8'h3;
initial mem[882] = 8'h3;
initial mem[883] = 8'h3;
initial mem[884] = 8'h3;
initial mem[885] = 8'h3;
initial mem[886] = 8'h3;
initial mem[887] = 8'h3;
initial mem[888] = 8'h3;
initial mem[889] = 8'h3;
initial mem[890] = 8'h3;
initial mem[891] = 8'h3;
initial mem[892] = 8'h3;
initial mem[893] = 8'h3;
initial mem[894] = 8'h3;
initial mem[895] = 8'h3;
initial mem[896] = 8'h3;
initial mem[897] = 8'h3;
initial mem[898] = 8'h3;
initial mem[899] = 8'h3;
initial mem[900] = 8'h3;
initial mem[901] = 8'h3;
initial mem[902] = 8'h3;
initial mem[903] = 8'h3;
initial mem[904] = 8'h3;
initial mem[905] = 8'h3;
initial mem[906] = 8'h3;
initial mem[907] = 8'h3;
initial mem[908] = 8'h3;
initial mem[909] = 8'h3;
initial mem[910] = 8'h3;
initial mem[911] = 8'h3;
initial mem[912] = 8'h3;
initial mem[913] = 8'h3;
initial mem[914] = 8'h3;
initial mem[915] = 8'h3;
initial mem[916] = 8'h3;
initial mem[917] = 8'h3;
initial mem[918] = 8'h3;
initial mem[919] = 8'h3;
initial mem[920] = 8'h3;
initial mem[921] = 8'h3;
initial mem[922] = 8'h3;
initial mem[923] = 8'h3;
initial mem[924] = 8'h3;
initial mem[925] = 8'h3;
initial mem[926] = 8'h3;
initial mem[927] = 8'h3;
initial mem[928] = 8'h3;
initial mem[929] = 8'h3;
initial mem[930] = 8'h3;
initial mem[931] = 8'h3;
initial mem[932] = 8'h3;
initial mem[933] = 8'h3;
initial mem[934] = 8'h3;
initial mem[935] = 8'h3;
initial mem[936] = 8'h3;
initial mem[937] = 8'h3;
initial mem[938] = 8'h3;
initial mem[939] = 8'h3;
initial mem[940] = 8'h3;
initial mem[941] = 8'h3;
initial mem[942] = 8'h3;
initial mem[943] = 8'h3;
initial mem[944] = 8'h3;
initial mem[945] = 8'h3;
initial mem[946] = 8'h3;
initial mem[947] = 8'h3;
initial mem[948] = 8'h3;
initial mem[949] = 8'h3;
initial mem[950] = 8'h3;
initial mem[951] = 8'h3;
initial mem[952] = 8'h3;
initial mem[953] = 8'h3;
initial mem[954] = 8'h3;
initial mem[955] = 8'h3;
initial mem[956] = 8'h3;
initial mem[957] = 8'h3;
initial mem[958] = 8'h3;
initial mem[959] = 8'h3;
initial mem[960] = 8'h3;
initial mem[961] = 8'h3;
initial mem[962] = 8'h3;
initial mem[963] = 8'h3;
initial mem[964] = 8'h3;
initial mem[965] = 8'h3;
initial mem[966] = 8'h3;
initial mem[967] = 8'h3;
initial mem[968] = 8'h3;
initial mem[969] = 8'h3;
initial mem[970] = 8'h3;
initial mem[971] = 8'h3;
initial mem[972] = 8'h3;
initial mem[973] = 8'h3;
initial mem[974] = 8'h3;
initial mem[975] = 8'h3;
initial mem[976] = 8'h3;
initial mem[977] = 8'h3;
initial mem[978] = 8'h3;
initial mem[979] = 8'h3;
initial mem[980] = 8'h3;
initial mem[981] = 8'h3;
initial mem[982] = 8'h3;
initial mem[983] = 8'h3;
initial mem[984] = 8'h3;
initial mem[985] = 8'h3;
initial mem[986] = 8'h3;
initial mem[987] = 8'h3;
initial mem[988] = 8'h3;
initial mem[989] = 8'h3;
initial mem[990] = 8'h3;
initial mem[991] = 8'h3;
initial mem[992] = 8'h3;
initial mem[993] = 8'h3;
initial mem[994] = 8'h3;
initial mem[995] = 8'h3;
initial mem[996] = 8'h3;
initial mem[997] = 8'h3;
initial mem[998] = 8'h3;
initial mem[999] = 8'h3;
initial mem[1000] = 8'h3;
initial mem[1001] = 8'h3;
initial mem[1002] = 8'h3;
initial mem[1003] = 8'h3;
initial mem[1004] = 8'h3;
initial mem[1005] = 8'h3;
initial mem[1006] = 8'h3;
initial mem[1007] = 8'h3;
initial mem[1008] = 8'h3;
initial mem[1009] = 8'h3;
initial mem[1010] = 8'h3;
initial mem[1011] = 8'h3;
initial mem[1012] = 8'h3;
initial mem[1013] = 8'h3;
initial mem[1014] = 8'h3;
initial mem[1015] = 8'h3;
initial mem[1016] = 8'h3;
initial mem[1017] = 8'h3;
initial mem[1018] = 8'h3;
initial mem[1019] = 8'h3;
initial mem[1020] = 8'h3;
initial mem[1021] = 8'h3;
initial mem[1022] = 8'h3;
initial mem[1023] = 8'h3;
always @(posedge clk) begin
	data <= mem[addr];
end
endmodule
